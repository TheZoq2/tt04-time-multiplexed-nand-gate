module \std::io::rising_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::rising_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::rising_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:3,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:4,14" *)
    logic _e_6;
    (* src = "<compiler dir>/stdlib/io.spade:4,5" *)
    logic _e_4;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_6 = !\sync2 ;
    assign _e_4 = \sync1  && _e_6;
    assign output__ = _e_4;
endmodule

module \std::io::falling_edge  (
        input clk_i,
        input sync1_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "std::io::falling_edge" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \std::io::falling_edge );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \sync1 ;
    assign \sync1  = sync1_i;
    (* src = "<compiler dir>/stdlib/io.spade:9,14" *)
    reg \sync2 ;
    (* src = "<compiler dir>/stdlib/io.spade:10,14" *)
    logic _e_14;
    (* src = "<compiler dir>/stdlib/io.spade:10,5" *)
    logic _e_12;
    always @(posedge \clk ) begin
        \sync2  <= \sync1 ;
    end
    assign _e_14 = !\sync1 ;
    assign _e_12 = \sync2  && _e_14;
    assign output__ = _e_12;
endmodule

module \tto4_tmng::main::regfile  (
        input clk_i,
        input[6:0] addr_i,
        input[8:0] write_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::main::regfile" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::main::regfile );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic[6:0] \addr ;
    assign \addr  = addr_i;
    logic[8:0] \write ;
    assign \write  = write_i;
    (* src = "src/main.spade:40,5" *)
    reg[6:0] \s1_addr ;
    (* src = "src/main.spade:40,5" *)
    reg[8:0] \s1_write ;
    (* src = "src/main.spade:40,5" *)
    reg[8:0] \s1_write_raw ;
    (* src = "src/main.spade:40,5" *)
    reg \s1_out ;
    logic[7:0] _e_62;
    logic[6:0] addr_n1;
    logic \b ;
    logic _e_3752;
    logic _e_3754;
    logic _e_3755;
    logic _e_3756;
    logic _e_3757;
    logic _e_65;
    (* src = "src/main.spade:33,33" *)
    logic[8:0] _e_64;
    logic _e_3759;
    logic _e_70;
    logic[6:0] _e_71;
    logic _e_72;
    (* src = "src/main.spade:34,22" *)
    logic[8:0] _e_69;
    (* src = "src/main.spade:32,25" *)
    logic[8:0] \write_raw ;
    (* src = "src/main.spade:37,63" *)
    logic[8:0] _e_76;
    (* src = "src/main.spade:37,38" *)
    logic[127:0] \mem ;
    (* src = "src/main.spade:39,19" *)
    logic \out ;
    logic[6:0] _e_3761;
    logic _e_3760;
    logic _e_86;
    logic[6:0] _e_3763;
    logic _e_3762;
    logic _e_88;
    logic _e_3764;
    (* src = "src/main.spade:41,9" *)
    logic _e_83;
    always @(posedge \clk ) begin
        \s1_addr  <= \addr ;
    end
    always @(posedge \clk ) begin
        \s1_write  <= \write ;
    end
    always @(posedge \clk ) begin
        \s1_write_raw  <= \write_raw ;
    end
    always @(posedge \clk ) begin
        \s1_out  <= \out ;
    end
    assign _e_62 = \write [7:0];
    assign addr_n1 = _e_62[7:1];
    assign \b  = _e_62[0];
    assign _e_3752 = \write [8] == 1'd0;
    assign _e_3754 = 1;
    assign _e_3755 = 1;
    assign _e_3756 = _e_3754 && _e_3755;
    assign _e_3757 = _e_3752 && _e_3756;
    assign _e_65 = 1;
    assign _e_64 = {_e_65, addr_n1, \b };
    assign _e_3759 = \write [8] == 1'd1;
    assign _e_70 = 0;
    assign _e_71 = 0;
    assign _e_72 = 0;
    assign _e_69 = {_e_70, _e_71, _e_72};
    always_comb begin
        priority casez ({_e_3757, _e_3759})
            2'b1?: \write_raw  = _e_64;
            2'b01: \write_raw  = _e_69;
            2'b?: \write_raw  = 'x;
        endcase
    end
    assign _e_76 = {\write_raw };
    always @(posedge \clk ) begin
        if (_e_76[8]) begin
            \mem [_e_76[7:1]] <= _e_76[0];
        end
    end
    assign \out  = \mem [\addr ];
    assign _e_3761 = 0;
    assign _e_3760 = \s1_addr  == _e_3761;
    assign _e_86 = 0;
    assign _e_3763 = 1;
    assign _e_3762 = \s1_addr  == _e_3763;
    assign _e_88 = 1;
    assign _e_3764 = 1;
    always_comb begin
        priority casez ({_e_3760, _e_3762, _e_3764})
            3'b1??: _e_83 = _e_86;
            3'b01?: _e_83 = _e_88;
            3'b001: _e_83 = \s1_out ;
            3'b?: _e_83 = 'x;
        endcase
    end
    assign output__ = _e_83;
endmodule

module \tto4_tmng::main::decode_extra_control  (
        input clk_i,
        input mode_i,
        input[7:0] uio_in_i,
        output output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::main::decode_extra_control" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::main::decode_extra_control );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \mode ;
    assign \mode  = mode_i;
    logic[7:0] \uio_in ;
    assign \uio_in  = uio_in_i;
    logic[7:0] _e_102;
    (* src = "src/main.spade:55,63" *)
    logic[7:0] _e_100;
    logic[7:0] _e_103;
    (* src = "src/main.spade:55,63" *)
    logic _e_99;
    (* src = "src/main.spade:55,31" *)
    logic _e_94;
    (* src = "src/main.spade:55,14" *)
    reg \push_to_output ;
    (* src = "src/main.spade:57,5" *)
    logic _e_104;
    assign _e_102 = 1;
    assign _e_100 = \uio_in  & _e_102;
    assign _e_103 = 1;
    assign _e_99 = _e_100 == _e_103;
    assign _e_94 = \mode  ? \push_to_output  : _e_99;
    always @(posedge \clk ) begin
        \push_to_output  <= _e_94;
    end
    assign _e_104 = {\push_to_output };
    assign output__ = _e_104;
endmodule

module \tto4_tmng::main::output_fifo  (
        input clk_i,
        input[1:0] push_i,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::main::output_fifo" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::main::output_fifo );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic[1:0] \push ;
    assign \push  = push_i;
    logic \next ;
    logic _e_3766;
    logic _e_3767;
    logic _e_3768;
    logic[7:0] _e_116;
    (* src = "src/main.spade:64,23" *)
    logic[7:0] _e_114;
    logic[7:0] _e_120;
    logic[7:0] _e_122;
    (* src = "src/main.spade:64,38" *)
    logic[7:0] _e_117;
    (* src = "src/main.spade:64,23" *)
    logic[7:0] _e_113;
    logic _e_3770;
    (* src = "src/main.spade:63,24" *)
    logic[7:0] _e_109;
    (* src = "src/main.spade:63,14" *)
    reg[7:0] \content ;
    assign \next  = \push [0:0];
    assign _e_3766 = \push [1] == 1'd0;
    assign _e_3767 = 1;
    assign _e_3768 = _e_3766 && _e_3767;
    assign _e_116 = 1;
    assign _e_114 = \content  << _e_116;
    assign _e_120 = 1;
    assign _e_122 = 0;
    assign _e_117 = \next  ? _e_120 : _e_122;
    assign _e_113 = _e_114 | _e_117;
    assign _e_3770 = \push [1] == 1'd1;
    always_comb begin
        priority casez ({_e_3768, _e_3770})
            2'b1?: _e_109 = _e_113;
            2'b01: _e_109 = \content ;
            2'b?: _e_109 = 'x;
        endcase
    end
    always @(posedge \clk ) begin
        \content  <= _e_109;
    end
    assign output__ = \content ;
endmodule

module \tto4_tmng::main::top_impl  (
        input clk_i,
        input[7:0] ui_in_i,
        input[7:0] uio_in_i,
        output[8:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::main::top_impl" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::main::top_impl );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic[7:0] \ui_in ;
    assign \ui_in  = ui_in_i;
    logic[7:0] \uio_in ;
    assign \uio_in  = uio_in_i;
    (* src = "src/main.spade:83,5" *)
    reg[7:0] \s1_ui_in ;
    (* src = "src/main.spade:83,5" *)
    reg[7:0] \s1_uio_in ;
    (* src = "src/main.spade:84,5" *)
    reg[7:0] \s2_ui_in ;
    (* src = "src/main.spade:84,5" *)
    reg[7:0] \s2_uio_in ;
    (* src = "src/main.spade:103,5" *)
    reg[7:0] \s3_ui_in ;
    (* src = "src/main.spade:103,5" *)
    reg[7:0] \s3_uio_in ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_mode ;
    (* src = "src/main.spade:103,5" *)
    reg[6:0] \s3_addr1 ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_commit_raw ;
    (* src = "src/main.spade:103,5" *)
    reg[6:0] \s3_addr2 ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_extra_control ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_commit_old ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_commit ;
    (* src = "src/main.spade:103,5" *)
    reg \s3_wb ;
    (* src = "src/main.spade:103,5" *)
    reg[6:0] \s3_wb_addr ;
    (* src = "src/main.spade:103,5" *)
    reg[8:0] \s3_write ;
    logic[7:0] _e_132;
    (* src = "src/main.spade:85,32" *)
    logic[7:0] _e_130;
    logic[7:0] _e_133;
    (* src = "src/main.spade:85,32" *)
    logic[7:0] _e_129;
    logic[7:0] _e_134;
    (* src = "src/main.spade:85,32" *)
    logic _e_128;
    (* src = "src/main.spade:85,55" *)
    logic[6:0] _e_135;
    (* src = "src/main.spade:85,32" *)
    logic[7:0] _e_139;
    logic \mode ;
    logic[6:0] \addr1 ;
    logic[7:0] _e_145;
    (* src = "src/main.spade:86,38" *)
    logic[7:0] _e_143;
    logic[7:0] _e_146;
    (* src = "src/main.spade:86,38" *)
    logic[7:0] _e_142;
    logic[7:0] _e_147;
    (* src = "src/main.spade:86,38" *)
    logic _e_141;
    (* src = "src/main.spade:86,62" *)
    logic[6:0] _e_148;
    (* src = "src/main.spade:86,38" *)
    logic[7:0] _e_152;
    logic \commit_raw ;
    logic[6:0] \addr2 ;
    (* src = "src/main.spade:88,29" *)
    logic \extra_control ;
    (* src = "src/main.spade:90,18" *)
    reg \commit_old ;
    (* src = "src/main.spade:91,36" *)
    logic _e_163;
    (* src = "src/main.spade:91,22" *)
    logic \commit ;
    (* src = "src/main.spade:93,13" *)
    logic \wb ;
    (* src = "src/main.spade:94,13" *)
    logic[6:0] \wb_addr ;
    (* src = "src/main.spade:95,24" *)
    logic _e_171;
    (* src = "src/main.spade:96,19" *)
    logic[7:0] _e_176;
    (* src = "src/main.spade:96,13" *)
    logic[8:0] _e_175;
    (* src = "src/main.spade:99,13" *)
    logic[8:0] _e_180;
    (* src = "src/main.spade:95,21" *)
    logic[8:0] \write ;
    (* src = "src/main.spade:102,23" *)
    logic \reg_out ;
    (* src = "src/main.spade:106,27" *)
    logic _e_190;
    (* src = "src/main.spade:106,24" *)
    logic _e_189;
    (* src = "src/main.spade:106,18" *)
    reg \opa ;
    (* src = "src/main.spade:107,13" *)
    logic \opb ;
    (* src = "src/main.spade:109,26" *)
    logic _e_199;
    (* src = "src/main.spade:109,24" *)
    logic \nand_out ;
    (* src = "src/main.spade:113,16" *)
    logic _e_207;
    (* src = "src/main.spade:113,16" *)
    logic _e_206;
    (* src = "src/main.spade:113,56" *)
    logic[1:0] _e_211;
    (* src = "src/main.spade:113,78" *)
    logic[1:0] _e_214;
    (* src = "src/main.spade:113,13" *)
    logic[1:0] _e_205;
    (* src = "src/main.spade:111,27" *)
    logic[7:0] \output_bits ;
    (* src = "src/main.spade:116,31" *)
    logic _e_218;
    (* src = "src/main.spade:116,18" *)
    reg \nand_snoop ;
    (* src = "src/main.spade:118,9" *)
    logic[8:0] _e_224;
    always @(posedge \clk ) begin
        \s1_ui_in  <= \ui_in ;
    end
    always @(posedge \clk ) begin
        \s1_uio_in  <= \uio_in ;
    end
    always @(posedge \clk ) begin
        \s2_ui_in  <= \s1_ui_in ;
    end
    always @(posedge \clk ) begin
        \s2_uio_in  <= \s1_uio_in ;
    end
    always @(posedge \clk ) begin
        \s3_ui_in  <= \s2_ui_in ;
    end
    always @(posedge \clk ) begin
        \s3_uio_in  <= \s2_uio_in ;
    end
    always @(posedge \clk ) begin
        \s3_mode  <= \mode ;
    end
    always @(posedge \clk ) begin
        \s3_addr1  <= \addr1 ;
    end
    always @(posedge \clk ) begin
        \s3_commit_raw  <= \commit_raw ;
    end
    always @(posedge \clk ) begin
        \s3_addr2  <= \addr2 ;
    end
    always @(posedge \clk ) begin
        \s3_extra_control  <= \extra_control ;
    end
    always @(posedge \clk ) begin
        \s3_commit_old  <= \commit_old ;
    end
    always @(posedge \clk ) begin
        \s3_commit  <= \commit ;
    end
    always @(posedge \clk ) begin
        \s3_wb  <= \wb ;
    end
    always @(posedge \clk ) begin
        \s3_wb_addr  <= \wb_addr ;
    end
    always @(posedge \clk ) begin
        \s3_write  <= \write ;
    end
    assign _e_132 = 7;
    assign _e_130 = \s2_ui_in  >> _e_132;
    assign _e_133 = 1;
    assign _e_129 = _e_130 & _e_133;
    assign _e_134 = 1;
    assign _e_128 = _e_129 == _e_134;
    assign _e_135 = \s2_ui_in [6:0];
    assign _e_139 = {_e_128, _e_135};
    assign \mode  = _e_139[7];
    assign \addr1  = _e_139[6:0];
    assign _e_145 = 7;
    assign _e_143 = \s2_uio_in  >> _e_145;
    assign _e_146 = 1;
    assign _e_142 = _e_143 & _e_146;
    assign _e_147 = 1;
    assign _e_141 = _e_142 == _e_147;
    assign _e_148 = \s2_uio_in [6:0];
    assign _e_152 = {_e_141, _e_148};
    assign \commit_raw  = _e_152[7];
    assign \addr2  = _e_152[6:0];
    (* src = "src/main.spade:88,29" *)
    \tto4_tmng::main::decode_extra_control  decode_extra_control_0(\clk , \mode , \s2_uio_in , \extra_control );
    always @(posedge \clk ) begin
        \commit_old  <= \commit_raw ;
    end
    assign _e_163 = !\commit_old ;
    assign \commit  = \commit_raw  && _e_163;
    assign \wb  = \nand_out ;
    assign \wb_addr  = \s3_addr2 ;
    assign _e_171 = \s3_mode  && \s3_commit ;
    assign _e_176 = {\wb_addr , \wb };
    assign _e_175 = {1'd0, _e_176};
    assign _e_180 = {1'd1, 8'bX};
    assign \write  = _e_171 ? _e_175 : _e_180;
    (* src = "src/main.spade:102,23" *)
    \tto4_tmng::main::regfile  regfile_0(\clk , \addr1 , \write , \reg_out );
    assign _e_190 = !\s3_mode ;
    assign _e_189 = _e_190 ? \reg_out  : \opa ;
    always @(posedge \clk ) begin
        \opa  <= _e_189;
    end
    assign \opb  = \reg_out ;
    assign _e_199 = \opa  && \opb ;
    assign \nand_out  = !_e_199;
    assign _e_207 = \s3_extra_control ;
    assign _e_206 = _e_207 && \s3_commit ;
    assign _e_211 = {1'd0, \nand_out };
    assign _e_214 = {1'd1, 1'bX};
    assign _e_205 = _e_206 ? _e_211 : _e_214;
    (* src = "src/main.spade:111,27" *)
    \tto4_tmng::main::output_fifo  output_fifo_0(\clk , _e_205, \output_bits );
    assign _e_218 = \s3_commit  ? \nand_out  : \nand_snoop ;
    always @(posedge \clk ) begin
        \nand_snoop  <= _e_218;
    end
    assign _e_224 = {\output_bits , \nand_out };
    assign output__ = _e_224;
endmodule

module tt_um_thezoq2_tmng (
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input clk,
        input ena,
        input rst_n
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tt_um_thezoq2_tmng" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, tt_um_thezoq2_tmng);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    logic[7:0] _e_229;
    logic[7:0] _e_231;
    (* src = "src/main.spade:148,15" *)
    logic[8:0] \out ;
    (* src = "src/main.spade:150,18" *)
    logic[7:0] _e_238;
    assign _e_229 = 0;
    assign \uio_out_mut  = _e_229;
    assign _e_231 = 0;
    assign \uio_oe_mut  = _e_231;
    (* src = "src/main.spade:148,15" *)
    \tto4_tmng::main::top_impl  top_impl_0(\clk , \ui_in , \uio_in , \out );
    assign _e_238 = \out [8:1];
    assign \uo_out_mut  = _e_238;
endmodule

module \tto4_tmng::main::impl_harness  (
        input[7:0] ui_in,
        input[7:0] uio_in,
        output[7:0] uio_out,
        output[7:0] uio_oe,
        input clk,
        input ena,
        input rst_n,
        output[7:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::main::impl_harness" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::main::impl_harness );
        end
    end
    `endif
    logic[7:0] \uio_out_mut ;
    assign uio_out = \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    assign uio_oe = \uio_oe_mut ;
    logic[7:0] \uo_out_mut ;
    (* src = "src/main.spade:168,13" *)
    logic[7:0] _e_253;
    
    (* src = "src/main.spade:168,13" *)
    tt_um_thezoq2_tmng tt_um_thezoq2_tmng_0(\ui_in , \uo_out_mut , \uio_in , \uio_out_mut , \uio_oe_mut , \clk , \ena , \rst_n );
    assign _e_253 = \uo_out_mut ;
    assign output__ = _e_253;
endmodule

module top_fpgatest (
        input[7:0] ui_in,
        output[7:0] uo_out,
        input[7:0] uio_in,
        input clk,
        output[7:0] ui_in_drive,
        output[7:0] uio_in_drive,
        output[7:0] pmod7
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "top_fpgatest" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, top_fpgatest);
        end
    end
    `endif
    logic[7:0] \uo_out_mut ;
    assign uo_out = \uo_out_mut ;
    logic[7:0] \ui_in_drive_mut ;
    assign ui_in_drive = \ui_in_drive_mut ;
    logic[7:0] \uio_in_drive_mut ;
    assign uio_in_drive = \uio_in_drive_mut ;
    logic[7:0] \pmod7_mut ;
    assign pmod7 = \pmod7_mut ;
    logic[9:0] _e_258;
    logic[9:0] _e_262;
    (* src = "src/fpgatest.spade:86,50" *)
    logic _e_260;
    logic[9:0] _e_267;
    (* src = "src/fpgatest.spade:86,72" *)
    logic[10:0] _e_265;
    (* src = "src/fpgatest.spade:86,66" *)
    logic[9:0] _e_264;
    (* src = "src/fpgatest.spade:86,47" *)
    logic[9:0] _e_259;
    (* src = "src/fpgatest.spade:86,14" *)
    reg[9:0] \rst_count ;
    logic[9:0] _e_272;
    (* src = "src/fpgatest.spade:87,15" *)
    logic \rst ;
    logic[7:0] \uio_out_mut ;
    logic[7:0] \uio_oe_mut ;
    logic _e_285;
    (* src = "src/fpgatest.spade:103,16" *)
    logic _e_286;
    (* src = "src/fpgatest.spade:95,13" *)
    (* src = "src/fpgatest.spade:106,22" *)
    logic[15:0] \driver_out ;
    (* src = "src/fpgatest.spade:107,23" *)
    logic[7:0] _e_294;
    (* src = "src/fpgatest.spade:108,24" *)
    logic[7:0] _e_297;
    logic[7:0] _e_300;
    assign _e_258 = 5;
    assign _e_262 = 0;
    assign _e_260 = \rst_count  != _e_262;
    assign _e_267 = 1;
    assign _e_265 = $signed(\rst_count ) - $signed(_e_267);
    assign _e_264 = _e_265[9:0];
    assign _e_259 = _e_260 ? _e_264 : \rst_count ;
    initial begin
        \rst_count  = 'b0000000101;
    end
    always @(posedge \clk ) begin
        \rst_count  <= _e_259;
    end
    assign _e_272 = 0;
    assign \rst  = \rst_count  != _e_272;
    
    
    assign _e_285 = 1;
    assign _e_286 = !\rst ;
    (* src = "src/fpgatest.spade:95,13" *)
    tt_um_thezoq2_tmng tt_um_thezoq2_tmng_0(\ui_in , \uo_out_mut , \uio_in , \uio_out_mut , \uio_oe_mut , \clk , _e_285, _e_286);
    (* src = "src/fpgatest.spade:106,22" *)
    \tto4_tmng::generated_driver::simple_test_driver  simple_test_driver_0(\clk , \rst , \driver_out );
    assign _e_294 = \driver_out [15:8];
    assign \ui_in_drive_mut  = _e_294;
    assign _e_297 = \driver_out [7:0];
    assign \uio_in_drive_mut  = _e_297;
    assign _e_300 = \uo_out_mut ;
    assign \pmod7_mut  = _e_300;
endmodule

module \tto4_tmng::generated_driver::simple_test_driver  (
        input clk_i,
        input rst_i,
        output[15:0] output__
    );
    `ifdef COCOTB_SIM
    string __top_module;
    string __vcd_file;
    initial begin
        if ($value$plusargs("TOP_MODULE=%s", __top_module) && __top_module == "tto4_tmng::generated_driver::simple_test_driver" && $value$plusargs("VCD_FILENAME=%s", __vcd_file)) begin
            $dumpfile (__vcd_file);
            $dumpvars (0, \tto4_tmng::generated_driver::simple_test_driver );
        end
    end
    `endif
    logic \clk ;
    assign \clk  = clk_i;
    logic \rst ;
    assign \rst  = rst_i;
    (* src = "src/generated_driver.spade:1161,5" *)
    reg \s1_rst ;
    (* src = "src/generated_driver.spade:1161,5" *)
    reg[47:0] \s1_state ;
    (* src = "src/generated_driver.spade:1161,5" *)
    reg[14:0] \s1_read_idx ;
    (* src = "src/generated_driver.spade:1161,5" *)
    reg[15:0] \s1_mem_out ;
    logic[31:0] _e_307;
    (* src = "src/generated_driver.spade:15,35" *)
    logic[47:0] _e_306;
    logic[31:0] _e_310;
    logic _e_3772;
    logic[31:0] _e_3774;
    logic _e_3773;
    logic _e_3775;
    logic[14:0] _e_313;
    logic[31:0] _e_314;
    (* src = "src/generated_driver.spade:16,41" *)
    logic[47:0] _e_312;
    logic[31:0] \duration ;
    logic _e_3777;
    logic _e_3778;
    logic _e_3779;
    logic[31:0] _e_321;
    (* src = "src/generated_driver.spade:17,56" *)
    logic[32:0] _e_319;
    (* src = "src/generated_driver.spade:17,50" *)
    logic[31:0] _e_318;
    (* src = "src/generated_driver.spade:17,38" *)
    logic[47:0] _e_317;
    logic[14:0] _e_322;
    logic[31:0] _e_323;
    logic _e_3781;
    logic[14:0] _e_3783;
    logic _e_3782;
    logic[31:0] _e_3785;
    logic _e_3784;
    logic _e_3786;
    logic _e_3787;
    logic[31:0] _e_327;
    (* src = "src/generated_driver.spade:19,17" *)
    logic[47:0] _e_326;
    logic[14:0] \idx ;
    logic[31:0] _e_329;
    logic _e_3789;
    logic _e_3790;
    logic[31:0] _e_3792;
    logic _e_3791;
    logic _e_3793;
    logic _e_3794;
    logic[14:0] _e_336;
    (* src = "src/generated_driver.spade:22,34" *)
    logic[15:0] _e_334;
    (* src = "src/generated_driver.spade:22,28" *)
    logic[14:0] _e_333;
    logic[31:0] _e_337;
    (* src = "src/generated_driver.spade:22,17" *)
    logic[47:0] _e_332;
    logic[14:0] idx_n1;
    logic[31:0] duration_n1;
    logic _e_3796;
    logic _e_3797;
    logic _e_3798;
    logic _e_3799;
    logic _e_3800;
    (* src = "src/generated_driver.spade:25,28" *)
    logic[14:0] _e_343;
    logic[31:0] _e_348;
    (* src = "src/generated_driver.spade:25,46" *)
    logic[32:0] _e_346;
    (* src = "src/generated_driver.spade:25,40" *)
    logic[31:0] _e_345;
    (* src = "src/generated_driver.spade:25,17" *)
    logic[47:0] _e_342;
    (* src = "src/generated_driver.spade:15,53" *)
    logic[47:0] _e_308;
    (* src = "src/generated_driver.spade:15,18" *)
    reg[47:0] \state ;
    logic[14:0] idx_n2;
    logic[31:0] \_ ;
    logic _e_3802;
    logic _e_3803;
    logic _e_3804;
    logic _e_3805;
    logic _e_3806;
    logic[31:0] __n1;
    logic _e_3808;
    logic _e_3809;
    logic _e_3810;
    logic[14:0] _e_357;
    (* src = "src/generated_driver.spade:29,24" *)
    logic[14:0] \read_idx ;
    (* src = "src/generated_driver.spade:34,54" *)
    logic[7:0] _e_364;
    logic[7:0] _e_365;
    (* src = "src/generated_driver.spade:34,60" *)
    logic[15:0] _e_363;
    logic[7:0] _e_367;
    logic[7:0] _e_368;
    (* src = "src/generated_driver.spade:35,2" *)
    logic[15:0] _e_366;
    logic[7:0] _e_370;
    logic[7:0] _e_371;
    (* src = "src/generated_driver.spade:36,2" *)
    logic[15:0] _e_369;
    logic[7:0] _e_373;
    logic[7:0] _e_374;
    (* src = "src/generated_driver.spade:37,2" *)
    logic[15:0] _e_372;
    logic[7:0] _e_376;
    logic[7:0] _e_377;
    (* src = "src/generated_driver.spade:38,2" *)
    logic[15:0] _e_375;
    logic[7:0] _e_379;
    logic[7:0] _e_380;
    (* src = "src/generated_driver.spade:39,2" *)
    logic[15:0] _e_378;
    logic[7:0] _e_382;
    logic[7:0] _e_383;
    (* src = "src/generated_driver.spade:40,2" *)
    logic[15:0] _e_381;
    logic[7:0] _e_385;
    logic[7:0] _e_386;
    (* src = "src/generated_driver.spade:41,2" *)
    logic[15:0] _e_384;
    logic[7:0] _e_388;
    logic[7:0] _e_389;
    (* src = "src/generated_driver.spade:42,2" *)
    logic[15:0] _e_387;
    logic[7:0] _e_391;
    logic[7:0] _e_392;
    (* src = "src/generated_driver.spade:43,2" *)
    logic[15:0] _e_390;
    logic[7:0] _e_394;
    logic[7:0] _e_395;
    (* src = "src/generated_driver.spade:44,2" *)
    logic[15:0] _e_393;
    logic[7:0] _e_397;
    logic[7:0] _e_398;
    (* src = "src/generated_driver.spade:45,2" *)
    logic[15:0] _e_396;
    logic[7:0] _e_400;
    logic[7:0] _e_401;
    (* src = "src/generated_driver.spade:46,2" *)
    logic[15:0] _e_399;
    logic[7:0] _e_403;
    logic[7:0] _e_404;
    (* src = "src/generated_driver.spade:47,2" *)
    logic[15:0] _e_402;
    logic[7:0] _e_406;
    logic[7:0] _e_407;
    (* src = "src/generated_driver.spade:48,2" *)
    logic[15:0] _e_405;
    logic[7:0] _e_409;
    logic[7:0] _e_410;
    (* src = "src/generated_driver.spade:49,2" *)
    logic[15:0] _e_408;
    logic[7:0] _e_412;
    logic[7:0] _e_413;
    (* src = "src/generated_driver.spade:50,2" *)
    logic[15:0] _e_411;
    logic[7:0] _e_415;
    logic[7:0] _e_416;
    (* src = "src/generated_driver.spade:51,2" *)
    logic[15:0] _e_414;
    logic[7:0] _e_418;
    logic[7:0] _e_419;
    (* src = "src/generated_driver.spade:52,2" *)
    logic[15:0] _e_417;
    logic[7:0] _e_421;
    logic[7:0] _e_422;
    (* src = "src/generated_driver.spade:53,2" *)
    logic[15:0] _e_420;
    logic[7:0] _e_424;
    logic[7:0] _e_425;
    (* src = "src/generated_driver.spade:54,2" *)
    logic[15:0] _e_423;
    logic[7:0] _e_427;
    logic[7:0] _e_428;
    (* src = "src/generated_driver.spade:55,2" *)
    logic[15:0] _e_426;
    logic[7:0] _e_430;
    logic[7:0] _e_431;
    (* src = "src/generated_driver.spade:56,2" *)
    logic[15:0] _e_429;
    logic[7:0] _e_433;
    logic[7:0] _e_434;
    (* src = "src/generated_driver.spade:57,2" *)
    logic[15:0] _e_432;
    logic[7:0] _e_436;
    logic[7:0] _e_437;
    (* src = "src/generated_driver.spade:58,2" *)
    logic[15:0] _e_435;
    logic[7:0] _e_439;
    logic[7:0] _e_440;
    (* src = "src/generated_driver.spade:59,2" *)
    logic[15:0] _e_438;
    logic[7:0] _e_442;
    logic[7:0] _e_443;
    (* src = "src/generated_driver.spade:60,2" *)
    logic[15:0] _e_441;
    logic[7:0] _e_445;
    logic[7:0] _e_446;
    (* src = "src/generated_driver.spade:61,2" *)
    logic[15:0] _e_444;
    logic[7:0] _e_448;
    logic[7:0] _e_449;
    (* src = "src/generated_driver.spade:62,2" *)
    logic[15:0] _e_447;
    logic[7:0] _e_451;
    logic[7:0] _e_452;
    (* src = "src/generated_driver.spade:63,2" *)
    logic[15:0] _e_450;
    logic[7:0] _e_454;
    logic[7:0] _e_455;
    (* src = "src/generated_driver.spade:64,2" *)
    logic[15:0] _e_453;
    logic[7:0] _e_457;
    logic[7:0] _e_458;
    (* src = "src/generated_driver.spade:65,2" *)
    logic[15:0] _e_456;
    logic[7:0] _e_460;
    logic[7:0] _e_461;
    (* src = "src/generated_driver.spade:66,2" *)
    logic[15:0] _e_459;
    logic[7:0] _e_463;
    logic[7:0] _e_464;
    (* src = "src/generated_driver.spade:67,2" *)
    logic[15:0] _e_462;
    logic[7:0] _e_466;
    logic[7:0] _e_467;
    (* src = "src/generated_driver.spade:68,2" *)
    logic[15:0] _e_465;
    logic[7:0] _e_469;
    logic[7:0] _e_470;
    (* src = "src/generated_driver.spade:69,2" *)
    logic[15:0] _e_468;
    logic[7:0] _e_472;
    logic[7:0] _e_473;
    (* src = "src/generated_driver.spade:70,2" *)
    logic[15:0] _e_471;
    logic[7:0] _e_475;
    logic[7:0] _e_476;
    (* src = "src/generated_driver.spade:71,2" *)
    logic[15:0] _e_474;
    logic[7:0] _e_478;
    logic[7:0] _e_479;
    (* src = "src/generated_driver.spade:72,2" *)
    logic[15:0] _e_477;
    logic[7:0] _e_481;
    logic[7:0] _e_482;
    (* src = "src/generated_driver.spade:73,2" *)
    logic[15:0] _e_480;
    logic[7:0] _e_484;
    logic[7:0] _e_485;
    (* src = "src/generated_driver.spade:74,2" *)
    logic[15:0] _e_483;
    logic[7:0] _e_487;
    logic[7:0] _e_488;
    (* src = "src/generated_driver.spade:75,2" *)
    logic[15:0] _e_486;
    logic[7:0] _e_490;
    logic[7:0] _e_491;
    (* src = "src/generated_driver.spade:76,2" *)
    logic[15:0] _e_489;
    logic[7:0] _e_493;
    logic[7:0] _e_494;
    (* src = "src/generated_driver.spade:77,2" *)
    logic[15:0] _e_492;
    logic[7:0] _e_496;
    logic[7:0] _e_497;
    (* src = "src/generated_driver.spade:78,2" *)
    logic[15:0] _e_495;
    logic[7:0] _e_499;
    logic[7:0] _e_500;
    (* src = "src/generated_driver.spade:79,2" *)
    logic[15:0] _e_498;
    logic[7:0] _e_502;
    logic[7:0] _e_503;
    (* src = "src/generated_driver.spade:80,2" *)
    logic[15:0] _e_501;
    logic[7:0] _e_505;
    logic[7:0] _e_506;
    (* src = "src/generated_driver.spade:81,2" *)
    logic[15:0] _e_504;
    logic[7:0] _e_508;
    logic[7:0] _e_509;
    (* src = "src/generated_driver.spade:82,2" *)
    logic[15:0] _e_507;
    logic[7:0] _e_511;
    logic[7:0] _e_512;
    (* src = "src/generated_driver.spade:83,2" *)
    logic[15:0] _e_510;
    logic[7:0] _e_514;
    logic[7:0] _e_515;
    (* src = "src/generated_driver.spade:84,2" *)
    logic[15:0] _e_513;
    logic[7:0] _e_517;
    logic[7:0] _e_518;
    (* src = "src/generated_driver.spade:85,2" *)
    logic[15:0] _e_516;
    logic[7:0] _e_520;
    logic[7:0] _e_521;
    (* src = "src/generated_driver.spade:86,2" *)
    logic[15:0] _e_519;
    logic[7:0] _e_523;
    logic[7:0] _e_524;
    (* src = "src/generated_driver.spade:87,2" *)
    logic[15:0] _e_522;
    logic[7:0] _e_526;
    logic[7:0] _e_527;
    (* src = "src/generated_driver.spade:88,2" *)
    logic[15:0] _e_525;
    logic[7:0] _e_529;
    logic[7:0] _e_530;
    (* src = "src/generated_driver.spade:89,2" *)
    logic[15:0] _e_528;
    logic[7:0] _e_532;
    logic[7:0] _e_533;
    (* src = "src/generated_driver.spade:90,2" *)
    logic[15:0] _e_531;
    logic[7:0] _e_535;
    logic[7:0] _e_536;
    (* src = "src/generated_driver.spade:91,2" *)
    logic[15:0] _e_534;
    logic[7:0] _e_538;
    logic[7:0] _e_539;
    (* src = "src/generated_driver.spade:92,2" *)
    logic[15:0] _e_537;
    logic[7:0] _e_541;
    logic[7:0] _e_542;
    (* src = "src/generated_driver.spade:93,2" *)
    logic[15:0] _e_540;
    logic[7:0] _e_544;
    logic[7:0] _e_545;
    (* src = "src/generated_driver.spade:94,2" *)
    logic[15:0] _e_543;
    logic[7:0] _e_547;
    logic[7:0] _e_548;
    (* src = "src/generated_driver.spade:95,2" *)
    logic[15:0] _e_546;
    logic[7:0] _e_550;
    logic[7:0] _e_551;
    (* src = "src/generated_driver.spade:96,2" *)
    logic[15:0] _e_549;
    logic[7:0] _e_553;
    logic[7:0] _e_554;
    (* src = "src/generated_driver.spade:97,2" *)
    logic[15:0] _e_552;
    logic[7:0] _e_556;
    logic[7:0] _e_557;
    (* src = "src/generated_driver.spade:98,2" *)
    logic[15:0] _e_555;
    logic[7:0] _e_559;
    logic[7:0] _e_560;
    (* src = "src/generated_driver.spade:99,2" *)
    logic[15:0] _e_558;
    logic[7:0] _e_562;
    logic[7:0] _e_563;
    (* src = "src/generated_driver.spade:100,2" *)
    logic[15:0] _e_561;
    logic[7:0] _e_565;
    logic[7:0] _e_566;
    (* src = "src/generated_driver.spade:101,2" *)
    logic[15:0] _e_564;
    logic[7:0] _e_568;
    logic[7:0] _e_569;
    (* src = "src/generated_driver.spade:102,2" *)
    logic[15:0] _e_567;
    logic[7:0] _e_571;
    logic[7:0] _e_572;
    (* src = "src/generated_driver.spade:103,2" *)
    logic[15:0] _e_570;
    logic[7:0] _e_574;
    logic[7:0] _e_575;
    (* src = "src/generated_driver.spade:104,2" *)
    logic[15:0] _e_573;
    logic[7:0] _e_577;
    logic[7:0] _e_578;
    (* src = "src/generated_driver.spade:105,2" *)
    logic[15:0] _e_576;
    logic[7:0] _e_580;
    logic[7:0] _e_581;
    (* src = "src/generated_driver.spade:106,2" *)
    logic[15:0] _e_579;
    logic[7:0] _e_583;
    logic[7:0] _e_584;
    (* src = "src/generated_driver.spade:107,2" *)
    logic[15:0] _e_582;
    logic[7:0] _e_586;
    logic[7:0] _e_587;
    (* src = "src/generated_driver.spade:108,2" *)
    logic[15:0] _e_585;
    logic[7:0] _e_589;
    logic[7:0] _e_590;
    (* src = "src/generated_driver.spade:109,2" *)
    logic[15:0] _e_588;
    logic[7:0] _e_592;
    logic[7:0] _e_593;
    (* src = "src/generated_driver.spade:110,2" *)
    logic[15:0] _e_591;
    logic[7:0] _e_595;
    logic[7:0] _e_596;
    (* src = "src/generated_driver.spade:111,2" *)
    logic[15:0] _e_594;
    logic[7:0] _e_598;
    logic[7:0] _e_599;
    (* src = "src/generated_driver.spade:112,2" *)
    logic[15:0] _e_597;
    logic[7:0] _e_601;
    logic[7:0] _e_602;
    (* src = "src/generated_driver.spade:113,2" *)
    logic[15:0] _e_600;
    logic[7:0] _e_604;
    logic[7:0] _e_605;
    (* src = "src/generated_driver.spade:114,2" *)
    logic[15:0] _e_603;
    logic[7:0] _e_607;
    logic[7:0] _e_608;
    (* src = "src/generated_driver.spade:115,2" *)
    logic[15:0] _e_606;
    logic[7:0] _e_610;
    logic[7:0] _e_611;
    (* src = "src/generated_driver.spade:116,2" *)
    logic[15:0] _e_609;
    logic[7:0] _e_613;
    logic[7:0] _e_614;
    (* src = "src/generated_driver.spade:117,2" *)
    logic[15:0] _e_612;
    logic[7:0] _e_616;
    logic[7:0] _e_617;
    (* src = "src/generated_driver.spade:118,2" *)
    logic[15:0] _e_615;
    logic[7:0] _e_619;
    logic[7:0] _e_620;
    (* src = "src/generated_driver.spade:119,2" *)
    logic[15:0] _e_618;
    logic[7:0] _e_622;
    logic[7:0] _e_623;
    (* src = "src/generated_driver.spade:120,2" *)
    logic[15:0] _e_621;
    logic[7:0] _e_625;
    logic[7:0] _e_626;
    (* src = "src/generated_driver.spade:121,2" *)
    logic[15:0] _e_624;
    logic[7:0] _e_628;
    logic[7:0] _e_629;
    (* src = "src/generated_driver.spade:122,2" *)
    logic[15:0] _e_627;
    logic[7:0] _e_631;
    logic[7:0] _e_632;
    (* src = "src/generated_driver.spade:123,2" *)
    logic[15:0] _e_630;
    logic[7:0] _e_634;
    logic[7:0] _e_635;
    (* src = "src/generated_driver.spade:124,2" *)
    logic[15:0] _e_633;
    logic[7:0] _e_637;
    logic[7:0] _e_638;
    (* src = "src/generated_driver.spade:125,2" *)
    logic[15:0] _e_636;
    logic[7:0] _e_640;
    logic[7:0] _e_641;
    (* src = "src/generated_driver.spade:126,2" *)
    logic[15:0] _e_639;
    logic[7:0] _e_643;
    logic[7:0] _e_644;
    (* src = "src/generated_driver.spade:127,2" *)
    logic[15:0] _e_642;
    logic[7:0] _e_646;
    logic[7:0] _e_647;
    (* src = "src/generated_driver.spade:128,2" *)
    logic[15:0] _e_645;
    logic[7:0] _e_649;
    logic[7:0] _e_650;
    (* src = "src/generated_driver.spade:129,2" *)
    logic[15:0] _e_648;
    logic[7:0] _e_652;
    logic[7:0] _e_653;
    (* src = "src/generated_driver.spade:130,2" *)
    logic[15:0] _e_651;
    logic[7:0] _e_655;
    logic[7:0] _e_656;
    (* src = "src/generated_driver.spade:131,2" *)
    logic[15:0] _e_654;
    logic[7:0] _e_658;
    logic[7:0] _e_659;
    (* src = "src/generated_driver.spade:132,2" *)
    logic[15:0] _e_657;
    logic[7:0] _e_661;
    logic[7:0] _e_662;
    (* src = "src/generated_driver.spade:133,2" *)
    logic[15:0] _e_660;
    logic[7:0] _e_664;
    logic[7:0] _e_665;
    (* src = "src/generated_driver.spade:134,2" *)
    logic[15:0] _e_663;
    logic[7:0] _e_667;
    logic[7:0] _e_668;
    (* src = "src/generated_driver.spade:135,2" *)
    logic[15:0] _e_666;
    logic[7:0] _e_670;
    logic[7:0] _e_671;
    (* src = "src/generated_driver.spade:136,2" *)
    logic[15:0] _e_669;
    logic[7:0] _e_673;
    logic[7:0] _e_674;
    (* src = "src/generated_driver.spade:137,2" *)
    logic[15:0] _e_672;
    logic[7:0] _e_676;
    logic[7:0] _e_677;
    (* src = "src/generated_driver.spade:138,2" *)
    logic[15:0] _e_675;
    logic[7:0] _e_679;
    logic[7:0] _e_680;
    (* src = "src/generated_driver.spade:139,2" *)
    logic[15:0] _e_678;
    logic[7:0] _e_682;
    logic[7:0] _e_683;
    (* src = "src/generated_driver.spade:140,2" *)
    logic[15:0] _e_681;
    logic[7:0] _e_685;
    logic[7:0] _e_686;
    (* src = "src/generated_driver.spade:141,2" *)
    logic[15:0] _e_684;
    logic[7:0] _e_688;
    logic[7:0] _e_689;
    (* src = "src/generated_driver.spade:142,2" *)
    logic[15:0] _e_687;
    logic[7:0] _e_691;
    logic[7:0] _e_692;
    (* src = "src/generated_driver.spade:143,2" *)
    logic[15:0] _e_690;
    logic[7:0] _e_694;
    logic[7:0] _e_695;
    (* src = "src/generated_driver.spade:144,2" *)
    logic[15:0] _e_693;
    logic[7:0] _e_697;
    logic[7:0] _e_698;
    (* src = "src/generated_driver.spade:145,2" *)
    logic[15:0] _e_696;
    logic[7:0] _e_700;
    logic[7:0] _e_701;
    (* src = "src/generated_driver.spade:146,2" *)
    logic[15:0] _e_699;
    logic[7:0] _e_703;
    logic[7:0] _e_704;
    (* src = "src/generated_driver.spade:147,2" *)
    logic[15:0] _e_702;
    logic[7:0] _e_706;
    logic[7:0] _e_707;
    (* src = "src/generated_driver.spade:148,2" *)
    logic[15:0] _e_705;
    logic[7:0] _e_709;
    logic[7:0] _e_710;
    (* src = "src/generated_driver.spade:149,2" *)
    logic[15:0] _e_708;
    logic[7:0] _e_712;
    logic[7:0] _e_713;
    (* src = "src/generated_driver.spade:150,2" *)
    logic[15:0] _e_711;
    logic[7:0] _e_715;
    logic[7:0] _e_716;
    (* src = "src/generated_driver.spade:151,2" *)
    logic[15:0] _e_714;
    logic[7:0] _e_718;
    logic[7:0] _e_719;
    (* src = "src/generated_driver.spade:152,2" *)
    logic[15:0] _e_717;
    logic[7:0] _e_721;
    logic[7:0] _e_722;
    (* src = "src/generated_driver.spade:153,2" *)
    logic[15:0] _e_720;
    logic[7:0] _e_724;
    logic[7:0] _e_725;
    (* src = "src/generated_driver.spade:154,2" *)
    logic[15:0] _e_723;
    logic[7:0] _e_727;
    logic[7:0] _e_728;
    (* src = "src/generated_driver.spade:155,2" *)
    logic[15:0] _e_726;
    logic[7:0] _e_730;
    logic[7:0] _e_731;
    (* src = "src/generated_driver.spade:156,2" *)
    logic[15:0] _e_729;
    logic[7:0] _e_733;
    logic[7:0] _e_734;
    (* src = "src/generated_driver.spade:157,2" *)
    logic[15:0] _e_732;
    logic[7:0] _e_736;
    logic[7:0] _e_737;
    (* src = "src/generated_driver.spade:158,2" *)
    logic[15:0] _e_735;
    logic[7:0] _e_739;
    logic[7:0] _e_740;
    (* src = "src/generated_driver.spade:159,2" *)
    logic[15:0] _e_738;
    logic[7:0] _e_742;
    logic[7:0] _e_743;
    (* src = "src/generated_driver.spade:160,2" *)
    logic[15:0] _e_741;
    logic[7:0] _e_745;
    logic[7:0] _e_746;
    (* src = "src/generated_driver.spade:161,2" *)
    logic[15:0] _e_744;
    logic[7:0] _e_748;
    logic[7:0] _e_749;
    (* src = "src/generated_driver.spade:162,2" *)
    logic[15:0] _e_747;
    logic[7:0] _e_751;
    logic[7:0] _e_752;
    (* src = "src/generated_driver.spade:163,2" *)
    logic[15:0] _e_750;
    logic[7:0] _e_754;
    logic[7:0] _e_755;
    (* src = "src/generated_driver.spade:164,2" *)
    logic[15:0] _e_753;
    logic[7:0] _e_757;
    logic[7:0] _e_758;
    (* src = "src/generated_driver.spade:165,2" *)
    logic[15:0] _e_756;
    logic[7:0] _e_760;
    logic[7:0] _e_761;
    (* src = "src/generated_driver.spade:166,2" *)
    logic[15:0] _e_759;
    logic[7:0] _e_763;
    logic[7:0] _e_764;
    (* src = "src/generated_driver.spade:167,2" *)
    logic[15:0] _e_762;
    logic[7:0] _e_766;
    logic[7:0] _e_767;
    (* src = "src/generated_driver.spade:168,2" *)
    logic[15:0] _e_765;
    logic[7:0] _e_769;
    logic[7:0] _e_770;
    (* src = "src/generated_driver.spade:169,2" *)
    logic[15:0] _e_768;
    logic[7:0] _e_772;
    logic[7:0] _e_773;
    (* src = "src/generated_driver.spade:170,2" *)
    logic[15:0] _e_771;
    logic[7:0] _e_775;
    logic[7:0] _e_776;
    (* src = "src/generated_driver.spade:171,2" *)
    logic[15:0] _e_774;
    logic[7:0] _e_778;
    logic[7:0] _e_779;
    (* src = "src/generated_driver.spade:172,2" *)
    logic[15:0] _e_777;
    logic[7:0] _e_781;
    logic[7:0] _e_782;
    (* src = "src/generated_driver.spade:173,2" *)
    logic[15:0] _e_780;
    logic[7:0] _e_784;
    logic[7:0] _e_785;
    (* src = "src/generated_driver.spade:174,2" *)
    logic[15:0] _e_783;
    logic[7:0] _e_787;
    logic[7:0] _e_788;
    (* src = "src/generated_driver.spade:175,2" *)
    logic[15:0] _e_786;
    logic[7:0] _e_790;
    logic[7:0] _e_791;
    (* src = "src/generated_driver.spade:176,2" *)
    logic[15:0] _e_789;
    logic[7:0] _e_793;
    logic[7:0] _e_794;
    (* src = "src/generated_driver.spade:177,2" *)
    logic[15:0] _e_792;
    logic[7:0] _e_796;
    logic[7:0] _e_797;
    (* src = "src/generated_driver.spade:178,2" *)
    logic[15:0] _e_795;
    logic[7:0] _e_799;
    logic[7:0] _e_800;
    (* src = "src/generated_driver.spade:179,2" *)
    logic[15:0] _e_798;
    logic[7:0] _e_802;
    logic[7:0] _e_803;
    (* src = "src/generated_driver.spade:180,2" *)
    logic[15:0] _e_801;
    logic[7:0] _e_805;
    logic[7:0] _e_806;
    (* src = "src/generated_driver.spade:181,2" *)
    logic[15:0] _e_804;
    logic[7:0] _e_808;
    logic[7:0] _e_809;
    (* src = "src/generated_driver.spade:182,2" *)
    logic[15:0] _e_807;
    logic[7:0] _e_811;
    logic[7:0] _e_812;
    (* src = "src/generated_driver.spade:183,2" *)
    logic[15:0] _e_810;
    logic[7:0] _e_814;
    logic[7:0] _e_815;
    (* src = "src/generated_driver.spade:184,2" *)
    logic[15:0] _e_813;
    logic[7:0] _e_817;
    logic[7:0] _e_818;
    (* src = "src/generated_driver.spade:185,2" *)
    logic[15:0] _e_816;
    logic[7:0] _e_820;
    logic[7:0] _e_821;
    (* src = "src/generated_driver.spade:186,2" *)
    logic[15:0] _e_819;
    logic[7:0] _e_823;
    logic[7:0] _e_824;
    (* src = "src/generated_driver.spade:187,2" *)
    logic[15:0] _e_822;
    logic[7:0] _e_826;
    logic[7:0] _e_827;
    (* src = "src/generated_driver.spade:188,2" *)
    logic[15:0] _e_825;
    logic[7:0] _e_829;
    logic[7:0] _e_830;
    (* src = "src/generated_driver.spade:189,2" *)
    logic[15:0] _e_828;
    logic[7:0] _e_832;
    logic[7:0] _e_833;
    (* src = "src/generated_driver.spade:190,2" *)
    logic[15:0] _e_831;
    logic[7:0] _e_835;
    logic[7:0] _e_836;
    (* src = "src/generated_driver.spade:191,2" *)
    logic[15:0] _e_834;
    logic[7:0] _e_838;
    logic[7:0] _e_839;
    (* src = "src/generated_driver.spade:192,2" *)
    logic[15:0] _e_837;
    logic[7:0] _e_841;
    logic[7:0] _e_842;
    (* src = "src/generated_driver.spade:193,2" *)
    logic[15:0] _e_840;
    logic[7:0] _e_844;
    logic[7:0] _e_845;
    (* src = "src/generated_driver.spade:194,2" *)
    logic[15:0] _e_843;
    logic[7:0] _e_847;
    logic[7:0] _e_848;
    (* src = "src/generated_driver.spade:195,2" *)
    logic[15:0] _e_846;
    logic[7:0] _e_850;
    logic[7:0] _e_851;
    (* src = "src/generated_driver.spade:196,2" *)
    logic[15:0] _e_849;
    logic[7:0] _e_853;
    logic[7:0] _e_854;
    (* src = "src/generated_driver.spade:197,2" *)
    logic[15:0] _e_852;
    logic[7:0] _e_856;
    logic[7:0] _e_857;
    (* src = "src/generated_driver.spade:198,2" *)
    logic[15:0] _e_855;
    logic[7:0] _e_859;
    logic[7:0] _e_860;
    (* src = "src/generated_driver.spade:199,2" *)
    logic[15:0] _e_858;
    logic[7:0] _e_862;
    logic[7:0] _e_863;
    (* src = "src/generated_driver.spade:200,2" *)
    logic[15:0] _e_861;
    logic[7:0] _e_865;
    logic[7:0] _e_866;
    (* src = "src/generated_driver.spade:201,2" *)
    logic[15:0] _e_864;
    logic[7:0] _e_868;
    logic[7:0] _e_869;
    (* src = "src/generated_driver.spade:202,2" *)
    logic[15:0] _e_867;
    logic[7:0] _e_871;
    logic[7:0] _e_872;
    (* src = "src/generated_driver.spade:203,2" *)
    logic[15:0] _e_870;
    logic[7:0] _e_874;
    logic[7:0] _e_875;
    (* src = "src/generated_driver.spade:204,2" *)
    logic[15:0] _e_873;
    logic[7:0] _e_877;
    logic[7:0] _e_878;
    (* src = "src/generated_driver.spade:205,2" *)
    logic[15:0] _e_876;
    logic[7:0] _e_880;
    logic[7:0] _e_881;
    (* src = "src/generated_driver.spade:206,2" *)
    logic[15:0] _e_879;
    logic[7:0] _e_883;
    logic[7:0] _e_884;
    (* src = "src/generated_driver.spade:207,2" *)
    logic[15:0] _e_882;
    logic[7:0] _e_886;
    logic[7:0] _e_887;
    (* src = "src/generated_driver.spade:208,2" *)
    logic[15:0] _e_885;
    logic[7:0] _e_889;
    logic[7:0] _e_890;
    (* src = "src/generated_driver.spade:209,2" *)
    logic[15:0] _e_888;
    logic[7:0] _e_892;
    logic[7:0] _e_893;
    (* src = "src/generated_driver.spade:210,2" *)
    logic[15:0] _e_891;
    logic[7:0] _e_895;
    logic[7:0] _e_896;
    (* src = "src/generated_driver.spade:211,2" *)
    logic[15:0] _e_894;
    logic[7:0] _e_898;
    logic[7:0] _e_899;
    (* src = "src/generated_driver.spade:212,2" *)
    logic[15:0] _e_897;
    logic[7:0] _e_901;
    logic[7:0] _e_902;
    (* src = "src/generated_driver.spade:213,2" *)
    logic[15:0] _e_900;
    logic[7:0] _e_904;
    logic[7:0] _e_905;
    (* src = "src/generated_driver.spade:214,2" *)
    logic[15:0] _e_903;
    logic[7:0] _e_907;
    logic[7:0] _e_908;
    (* src = "src/generated_driver.spade:215,2" *)
    logic[15:0] _e_906;
    logic[7:0] _e_910;
    logic[7:0] _e_911;
    (* src = "src/generated_driver.spade:216,2" *)
    logic[15:0] _e_909;
    logic[7:0] _e_913;
    logic[7:0] _e_914;
    (* src = "src/generated_driver.spade:217,2" *)
    logic[15:0] _e_912;
    logic[7:0] _e_916;
    logic[7:0] _e_917;
    (* src = "src/generated_driver.spade:218,2" *)
    logic[15:0] _e_915;
    logic[7:0] _e_919;
    logic[7:0] _e_920;
    (* src = "src/generated_driver.spade:219,2" *)
    logic[15:0] _e_918;
    logic[7:0] _e_922;
    logic[7:0] _e_923;
    (* src = "src/generated_driver.spade:220,2" *)
    logic[15:0] _e_921;
    logic[7:0] _e_925;
    logic[7:0] _e_926;
    (* src = "src/generated_driver.spade:221,2" *)
    logic[15:0] _e_924;
    logic[7:0] _e_928;
    logic[7:0] _e_929;
    (* src = "src/generated_driver.spade:222,2" *)
    logic[15:0] _e_927;
    logic[7:0] _e_931;
    logic[7:0] _e_932;
    (* src = "src/generated_driver.spade:223,2" *)
    logic[15:0] _e_930;
    logic[7:0] _e_934;
    logic[7:0] _e_935;
    (* src = "src/generated_driver.spade:224,2" *)
    logic[15:0] _e_933;
    logic[7:0] _e_937;
    logic[7:0] _e_938;
    (* src = "src/generated_driver.spade:225,2" *)
    logic[15:0] _e_936;
    logic[7:0] _e_940;
    logic[7:0] _e_941;
    (* src = "src/generated_driver.spade:226,2" *)
    logic[15:0] _e_939;
    logic[7:0] _e_943;
    logic[7:0] _e_944;
    (* src = "src/generated_driver.spade:227,2" *)
    logic[15:0] _e_942;
    logic[7:0] _e_946;
    logic[7:0] _e_947;
    (* src = "src/generated_driver.spade:228,2" *)
    logic[15:0] _e_945;
    logic[7:0] _e_949;
    logic[7:0] _e_950;
    (* src = "src/generated_driver.spade:229,2" *)
    logic[15:0] _e_948;
    logic[7:0] _e_952;
    logic[7:0] _e_953;
    (* src = "src/generated_driver.spade:230,2" *)
    logic[15:0] _e_951;
    logic[7:0] _e_955;
    logic[7:0] _e_956;
    (* src = "src/generated_driver.spade:231,2" *)
    logic[15:0] _e_954;
    logic[7:0] _e_958;
    logic[7:0] _e_959;
    (* src = "src/generated_driver.spade:232,2" *)
    logic[15:0] _e_957;
    logic[7:0] _e_961;
    logic[7:0] _e_962;
    (* src = "src/generated_driver.spade:233,2" *)
    logic[15:0] _e_960;
    logic[7:0] _e_964;
    logic[7:0] _e_965;
    (* src = "src/generated_driver.spade:234,2" *)
    logic[15:0] _e_963;
    logic[7:0] _e_967;
    logic[7:0] _e_968;
    (* src = "src/generated_driver.spade:235,2" *)
    logic[15:0] _e_966;
    logic[7:0] _e_970;
    logic[7:0] _e_971;
    (* src = "src/generated_driver.spade:236,2" *)
    logic[15:0] _e_969;
    logic[7:0] _e_973;
    logic[7:0] _e_974;
    (* src = "src/generated_driver.spade:237,2" *)
    logic[15:0] _e_972;
    logic[7:0] _e_976;
    logic[7:0] _e_977;
    (* src = "src/generated_driver.spade:238,2" *)
    logic[15:0] _e_975;
    logic[7:0] _e_979;
    logic[7:0] _e_980;
    (* src = "src/generated_driver.spade:239,2" *)
    logic[15:0] _e_978;
    logic[7:0] _e_982;
    logic[7:0] _e_983;
    (* src = "src/generated_driver.spade:240,2" *)
    logic[15:0] _e_981;
    logic[7:0] _e_985;
    logic[7:0] _e_986;
    (* src = "src/generated_driver.spade:241,2" *)
    logic[15:0] _e_984;
    logic[7:0] _e_988;
    logic[7:0] _e_989;
    (* src = "src/generated_driver.spade:242,2" *)
    logic[15:0] _e_987;
    logic[7:0] _e_991;
    logic[7:0] _e_992;
    (* src = "src/generated_driver.spade:243,2" *)
    logic[15:0] _e_990;
    logic[7:0] _e_994;
    logic[7:0] _e_995;
    (* src = "src/generated_driver.spade:244,2" *)
    logic[15:0] _e_993;
    logic[7:0] _e_997;
    logic[7:0] _e_998;
    (* src = "src/generated_driver.spade:245,2" *)
    logic[15:0] _e_996;
    logic[7:0] _e_1000;
    logic[7:0] _e_1001;
    (* src = "src/generated_driver.spade:246,2" *)
    logic[15:0] _e_999;
    logic[7:0] _e_1003;
    logic[7:0] _e_1004;
    (* src = "src/generated_driver.spade:247,2" *)
    logic[15:0] _e_1002;
    logic[7:0] _e_1006;
    logic[7:0] _e_1007;
    (* src = "src/generated_driver.spade:248,2" *)
    logic[15:0] _e_1005;
    logic[7:0] _e_1009;
    logic[7:0] _e_1010;
    (* src = "src/generated_driver.spade:249,2" *)
    logic[15:0] _e_1008;
    logic[7:0] _e_1012;
    logic[7:0] _e_1013;
    (* src = "src/generated_driver.spade:250,2" *)
    logic[15:0] _e_1011;
    logic[7:0] _e_1015;
    logic[7:0] _e_1016;
    (* src = "src/generated_driver.spade:251,2" *)
    logic[15:0] _e_1014;
    logic[7:0] _e_1018;
    logic[7:0] _e_1019;
    (* src = "src/generated_driver.spade:252,2" *)
    logic[15:0] _e_1017;
    logic[7:0] _e_1021;
    logic[7:0] _e_1022;
    (* src = "src/generated_driver.spade:253,2" *)
    logic[15:0] _e_1020;
    logic[7:0] _e_1024;
    logic[7:0] _e_1025;
    (* src = "src/generated_driver.spade:254,2" *)
    logic[15:0] _e_1023;
    logic[7:0] _e_1027;
    logic[7:0] _e_1028;
    (* src = "src/generated_driver.spade:255,2" *)
    logic[15:0] _e_1026;
    logic[7:0] _e_1030;
    logic[7:0] _e_1031;
    (* src = "src/generated_driver.spade:256,2" *)
    logic[15:0] _e_1029;
    logic[7:0] _e_1033;
    logic[7:0] _e_1034;
    (* src = "src/generated_driver.spade:257,2" *)
    logic[15:0] _e_1032;
    logic[7:0] _e_1036;
    logic[7:0] _e_1037;
    (* src = "src/generated_driver.spade:258,2" *)
    logic[15:0] _e_1035;
    logic[7:0] _e_1039;
    logic[7:0] _e_1040;
    (* src = "src/generated_driver.spade:259,2" *)
    logic[15:0] _e_1038;
    logic[7:0] _e_1042;
    logic[7:0] _e_1043;
    (* src = "src/generated_driver.spade:260,2" *)
    logic[15:0] _e_1041;
    logic[7:0] _e_1045;
    logic[7:0] _e_1046;
    (* src = "src/generated_driver.spade:261,2" *)
    logic[15:0] _e_1044;
    logic[7:0] _e_1048;
    logic[7:0] _e_1049;
    (* src = "src/generated_driver.spade:262,2" *)
    logic[15:0] _e_1047;
    logic[7:0] _e_1051;
    logic[7:0] _e_1052;
    (* src = "src/generated_driver.spade:263,2" *)
    logic[15:0] _e_1050;
    logic[7:0] _e_1054;
    logic[7:0] _e_1055;
    (* src = "src/generated_driver.spade:264,2" *)
    logic[15:0] _e_1053;
    logic[7:0] _e_1057;
    logic[7:0] _e_1058;
    (* src = "src/generated_driver.spade:265,2" *)
    logic[15:0] _e_1056;
    logic[7:0] _e_1060;
    logic[7:0] _e_1061;
    (* src = "src/generated_driver.spade:266,2" *)
    logic[15:0] _e_1059;
    logic[7:0] _e_1063;
    logic[7:0] _e_1064;
    (* src = "src/generated_driver.spade:267,2" *)
    logic[15:0] _e_1062;
    logic[7:0] _e_1066;
    logic[7:0] _e_1067;
    (* src = "src/generated_driver.spade:268,2" *)
    logic[15:0] _e_1065;
    logic[7:0] _e_1069;
    logic[7:0] _e_1070;
    (* src = "src/generated_driver.spade:269,2" *)
    logic[15:0] _e_1068;
    logic[7:0] _e_1072;
    logic[7:0] _e_1073;
    (* src = "src/generated_driver.spade:270,2" *)
    logic[15:0] _e_1071;
    logic[7:0] _e_1075;
    logic[7:0] _e_1076;
    (* src = "src/generated_driver.spade:271,2" *)
    logic[15:0] _e_1074;
    logic[7:0] _e_1078;
    logic[7:0] _e_1079;
    (* src = "src/generated_driver.spade:272,2" *)
    logic[15:0] _e_1077;
    logic[7:0] _e_1081;
    logic[7:0] _e_1082;
    (* src = "src/generated_driver.spade:273,2" *)
    logic[15:0] _e_1080;
    logic[7:0] _e_1084;
    logic[7:0] _e_1085;
    (* src = "src/generated_driver.spade:274,2" *)
    logic[15:0] _e_1083;
    logic[7:0] _e_1087;
    logic[7:0] _e_1088;
    (* src = "src/generated_driver.spade:275,2" *)
    logic[15:0] _e_1086;
    logic[7:0] _e_1090;
    logic[7:0] _e_1091;
    (* src = "src/generated_driver.spade:276,2" *)
    logic[15:0] _e_1089;
    logic[7:0] _e_1093;
    logic[7:0] _e_1094;
    (* src = "src/generated_driver.spade:277,2" *)
    logic[15:0] _e_1092;
    logic[7:0] _e_1096;
    logic[7:0] _e_1097;
    (* src = "src/generated_driver.spade:278,2" *)
    logic[15:0] _e_1095;
    logic[7:0] _e_1099;
    logic[7:0] _e_1100;
    (* src = "src/generated_driver.spade:279,2" *)
    logic[15:0] _e_1098;
    logic[7:0] _e_1102;
    logic[7:0] _e_1103;
    (* src = "src/generated_driver.spade:280,2" *)
    logic[15:0] _e_1101;
    logic[7:0] _e_1105;
    logic[7:0] _e_1106;
    (* src = "src/generated_driver.spade:281,2" *)
    logic[15:0] _e_1104;
    logic[7:0] _e_1108;
    logic[7:0] _e_1109;
    (* src = "src/generated_driver.spade:282,2" *)
    logic[15:0] _e_1107;
    logic[7:0] _e_1111;
    logic[7:0] _e_1112;
    (* src = "src/generated_driver.spade:283,2" *)
    logic[15:0] _e_1110;
    logic[7:0] _e_1114;
    logic[7:0] _e_1115;
    (* src = "src/generated_driver.spade:284,2" *)
    logic[15:0] _e_1113;
    logic[7:0] _e_1117;
    logic[7:0] _e_1118;
    (* src = "src/generated_driver.spade:285,2" *)
    logic[15:0] _e_1116;
    logic[7:0] _e_1120;
    logic[7:0] _e_1121;
    (* src = "src/generated_driver.spade:286,2" *)
    logic[15:0] _e_1119;
    logic[7:0] _e_1123;
    logic[7:0] _e_1124;
    (* src = "src/generated_driver.spade:287,2" *)
    logic[15:0] _e_1122;
    logic[7:0] _e_1126;
    logic[7:0] _e_1127;
    (* src = "src/generated_driver.spade:288,2" *)
    logic[15:0] _e_1125;
    logic[7:0] _e_1129;
    logic[7:0] _e_1130;
    (* src = "src/generated_driver.spade:289,2" *)
    logic[15:0] _e_1128;
    logic[7:0] _e_1132;
    logic[7:0] _e_1133;
    (* src = "src/generated_driver.spade:290,2" *)
    logic[15:0] _e_1131;
    logic[7:0] _e_1135;
    logic[7:0] _e_1136;
    (* src = "src/generated_driver.spade:291,2" *)
    logic[15:0] _e_1134;
    logic[7:0] _e_1138;
    logic[7:0] _e_1139;
    (* src = "src/generated_driver.spade:292,2" *)
    logic[15:0] _e_1137;
    logic[7:0] _e_1141;
    logic[7:0] _e_1142;
    (* src = "src/generated_driver.spade:293,2" *)
    logic[15:0] _e_1140;
    logic[7:0] _e_1144;
    logic[7:0] _e_1145;
    (* src = "src/generated_driver.spade:294,2" *)
    logic[15:0] _e_1143;
    logic[7:0] _e_1147;
    logic[7:0] _e_1148;
    (* src = "src/generated_driver.spade:295,2" *)
    logic[15:0] _e_1146;
    logic[7:0] _e_1150;
    logic[7:0] _e_1151;
    (* src = "src/generated_driver.spade:296,2" *)
    logic[15:0] _e_1149;
    logic[7:0] _e_1153;
    logic[7:0] _e_1154;
    (* src = "src/generated_driver.spade:297,2" *)
    logic[15:0] _e_1152;
    logic[7:0] _e_1156;
    logic[7:0] _e_1157;
    (* src = "src/generated_driver.spade:298,2" *)
    logic[15:0] _e_1155;
    logic[7:0] _e_1159;
    logic[7:0] _e_1160;
    (* src = "src/generated_driver.spade:299,2" *)
    logic[15:0] _e_1158;
    logic[7:0] _e_1162;
    logic[7:0] _e_1163;
    (* src = "src/generated_driver.spade:300,2" *)
    logic[15:0] _e_1161;
    logic[7:0] _e_1165;
    logic[7:0] _e_1166;
    (* src = "src/generated_driver.spade:301,2" *)
    logic[15:0] _e_1164;
    logic[7:0] _e_1168;
    logic[7:0] _e_1169;
    (* src = "src/generated_driver.spade:302,2" *)
    logic[15:0] _e_1167;
    logic[7:0] _e_1171;
    logic[7:0] _e_1172;
    (* src = "src/generated_driver.spade:303,2" *)
    logic[15:0] _e_1170;
    logic[7:0] _e_1174;
    logic[7:0] _e_1175;
    (* src = "src/generated_driver.spade:304,2" *)
    logic[15:0] _e_1173;
    logic[7:0] _e_1177;
    logic[7:0] _e_1178;
    (* src = "src/generated_driver.spade:305,2" *)
    logic[15:0] _e_1176;
    logic[7:0] _e_1180;
    logic[7:0] _e_1181;
    (* src = "src/generated_driver.spade:306,2" *)
    logic[15:0] _e_1179;
    logic[7:0] _e_1183;
    logic[7:0] _e_1184;
    (* src = "src/generated_driver.spade:307,2" *)
    logic[15:0] _e_1182;
    logic[7:0] _e_1186;
    logic[7:0] _e_1187;
    (* src = "src/generated_driver.spade:308,2" *)
    logic[15:0] _e_1185;
    logic[7:0] _e_1189;
    logic[7:0] _e_1190;
    (* src = "src/generated_driver.spade:309,2" *)
    logic[15:0] _e_1188;
    logic[7:0] _e_1192;
    logic[7:0] _e_1193;
    (* src = "src/generated_driver.spade:310,2" *)
    logic[15:0] _e_1191;
    logic[7:0] _e_1195;
    logic[7:0] _e_1196;
    (* src = "src/generated_driver.spade:311,2" *)
    logic[15:0] _e_1194;
    logic[7:0] _e_1198;
    logic[7:0] _e_1199;
    (* src = "src/generated_driver.spade:312,2" *)
    logic[15:0] _e_1197;
    logic[7:0] _e_1201;
    logic[7:0] _e_1202;
    (* src = "src/generated_driver.spade:313,2" *)
    logic[15:0] _e_1200;
    logic[7:0] _e_1204;
    logic[7:0] _e_1205;
    (* src = "src/generated_driver.spade:314,2" *)
    logic[15:0] _e_1203;
    logic[7:0] _e_1207;
    logic[7:0] _e_1208;
    (* src = "src/generated_driver.spade:315,2" *)
    logic[15:0] _e_1206;
    logic[7:0] _e_1210;
    logic[7:0] _e_1211;
    (* src = "src/generated_driver.spade:316,2" *)
    logic[15:0] _e_1209;
    logic[7:0] _e_1213;
    logic[7:0] _e_1214;
    (* src = "src/generated_driver.spade:317,2" *)
    logic[15:0] _e_1212;
    logic[7:0] _e_1216;
    logic[7:0] _e_1217;
    (* src = "src/generated_driver.spade:318,2" *)
    logic[15:0] _e_1215;
    logic[7:0] _e_1219;
    logic[7:0] _e_1220;
    (* src = "src/generated_driver.spade:319,2" *)
    logic[15:0] _e_1218;
    logic[7:0] _e_1222;
    logic[7:0] _e_1223;
    (* src = "src/generated_driver.spade:320,2" *)
    logic[15:0] _e_1221;
    logic[7:0] _e_1225;
    logic[7:0] _e_1226;
    (* src = "src/generated_driver.spade:321,2" *)
    logic[15:0] _e_1224;
    logic[7:0] _e_1228;
    logic[7:0] _e_1229;
    (* src = "src/generated_driver.spade:322,2" *)
    logic[15:0] _e_1227;
    logic[7:0] _e_1231;
    logic[7:0] _e_1232;
    (* src = "src/generated_driver.spade:323,2" *)
    logic[15:0] _e_1230;
    logic[7:0] _e_1234;
    logic[7:0] _e_1235;
    (* src = "src/generated_driver.spade:324,2" *)
    logic[15:0] _e_1233;
    logic[7:0] _e_1237;
    logic[7:0] _e_1238;
    (* src = "src/generated_driver.spade:325,2" *)
    logic[15:0] _e_1236;
    logic[7:0] _e_1240;
    logic[7:0] _e_1241;
    (* src = "src/generated_driver.spade:326,2" *)
    logic[15:0] _e_1239;
    logic[7:0] _e_1243;
    logic[7:0] _e_1244;
    (* src = "src/generated_driver.spade:327,2" *)
    logic[15:0] _e_1242;
    logic[7:0] _e_1246;
    logic[7:0] _e_1247;
    (* src = "src/generated_driver.spade:328,2" *)
    logic[15:0] _e_1245;
    logic[7:0] _e_1249;
    logic[7:0] _e_1250;
    (* src = "src/generated_driver.spade:329,2" *)
    logic[15:0] _e_1248;
    logic[7:0] _e_1252;
    logic[7:0] _e_1253;
    (* src = "src/generated_driver.spade:330,2" *)
    logic[15:0] _e_1251;
    logic[7:0] _e_1255;
    logic[7:0] _e_1256;
    (* src = "src/generated_driver.spade:331,2" *)
    logic[15:0] _e_1254;
    logic[7:0] _e_1258;
    logic[7:0] _e_1259;
    (* src = "src/generated_driver.spade:332,2" *)
    logic[15:0] _e_1257;
    logic[7:0] _e_1261;
    logic[7:0] _e_1262;
    (* src = "src/generated_driver.spade:333,2" *)
    logic[15:0] _e_1260;
    logic[7:0] _e_1264;
    logic[7:0] _e_1265;
    (* src = "src/generated_driver.spade:334,2" *)
    logic[15:0] _e_1263;
    logic[7:0] _e_1267;
    logic[7:0] _e_1268;
    (* src = "src/generated_driver.spade:335,2" *)
    logic[15:0] _e_1266;
    logic[7:0] _e_1270;
    logic[7:0] _e_1271;
    (* src = "src/generated_driver.spade:336,2" *)
    logic[15:0] _e_1269;
    logic[7:0] _e_1273;
    logic[7:0] _e_1274;
    (* src = "src/generated_driver.spade:337,2" *)
    logic[15:0] _e_1272;
    logic[7:0] _e_1276;
    logic[7:0] _e_1277;
    (* src = "src/generated_driver.spade:338,2" *)
    logic[15:0] _e_1275;
    logic[7:0] _e_1279;
    logic[7:0] _e_1280;
    (* src = "src/generated_driver.spade:339,2" *)
    logic[15:0] _e_1278;
    logic[7:0] _e_1282;
    logic[7:0] _e_1283;
    (* src = "src/generated_driver.spade:340,2" *)
    logic[15:0] _e_1281;
    logic[7:0] _e_1285;
    logic[7:0] _e_1286;
    (* src = "src/generated_driver.spade:341,2" *)
    logic[15:0] _e_1284;
    logic[7:0] _e_1288;
    logic[7:0] _e_1289;
    (* src = "src/generated_driver.spade:342,2" *)
    logic[15:0] _e_1287;
    logic[7:0] _e_1291;
    logic[7:0] _e_1292;
    (* src = "src/generated_driver.spade:343,2" *)
    logic[15:0] _e_1290;
    logic[7:0] _e_1294;
    logic[7:0] _e_1295;
    (* src = "src/generated_driver.spade:344,2" *)
    logic[15:0] _e_1293;
    logic[7:0] _e_1297;
    logic[7:0] _e_1298;
    (* src = "src/generated_driver.spade:345,2" *)
    logic[15:0] _e_1296;
    logic[7:0] _e_1300;
    logic[7:0] _e_1301;
    (* src = "src/generated_driver.spade:346,2" *)
    logic[15:0] _e_1299;
    logic[7:0] _e_1303;
    logic[7:0] _e_1304;
    (* src = "src/generated_driver.spade:347,2" *)
    logic[15:0] _e_1302;
    logic[7:0] _e_1306;
    logic[7:0] _e_1307;
    (* src = "src/generated_driver.spade:348,2" *)
    logic[15:0] _e_1305;
    logic[7:0] _e_1309;
    logic[7:0] _e_1310;
    (* src = "src/generated_driver.spade:349,2" *)
    logic[15:0] _e_1308;
    logic[7:0] _e_1312;
    logic[7:0] _e_1313;
    (* src = "src/generated_driver.spade:350,2" *)
    logic[15:0] _e_1311;
    logic[7:0] _e_1315;
    logic[7:0] _e_1316;
    (* src = "src/generated_driver.spade:351,2" *)
    logic[15:0] _e_1314;
    logic[7:0] _e_1318;
    logic[7:0] _e_1319;
    (* src = "src/generated_driver.spade:352,2" *)
    logic[15:0] _e_1317;
    logic[7:0] _e_1321;
    logic[7:0] _e_1322;
    (* src = "src/generated_driver.spade:353,2" *)
    logic[15:0] _e_1320;
    logic[7:0] _e_1324;
    logic[7:0] _e_1325;
    (* src = "src/generated_driver.spade:354,2" *)
    logic[15:0] _e_1323;
    logic[7:0] _e_1327;
    logic[7:0] _e_1328;
    (* src = "src/generated_driver.spade:355,2" *)
    logic[15:0] _e_1326;
    logic[7:0] _e_1330;
    logic[7:0] _e_1331;
    (* src = "src/generated_driver.spade:356,2" *)
    logic[15:0] _e_1329;
    logic[7:0] _e_1333;
    logic[7:0] _e_1334;
    (* src = "src/generated_driver.spade:357,2" *)
    logic[15:0] _e_1332;
    logic[7:0] _e_1336;
    logic[7:0] _e_1337;
    (* src = "src/generated_driver.spade:358,2" *)
    logic[15:0] _e_1335;
    logic[7:0] _e_1339;
    logic[7:0] _e_1340;
    (* src = "src/generated_driver.spade:359,2" *)
    logic[15:0] _e_1338;
    logic[7:0] _e_1342;
    logic[7:0] _e_1343;
    (* src = "src/generated_driver.spade:360,2" *)
    logic[15:0] _e_1341;
    logic[7:0] _e_1345;
    logic[7:0] _e_1346;
    (* src = "src/generated_driver.spade:361,2" *)
    logic[15:0] _e_1344;
    logic[7:0] _e_1348;
    logic[7:0] _e_1349;
    (* src = "src/generated_driver.spade:362,2" *)
    logic[15:0] _e_1347;
    logic[7:0] _e_1351;
    logic[7:0] _e_1352;
    (* src = "src/generated_driver.spade:363,2" *)
    logic[15:0] _e_1350;
    logic[7:0] _e_1354;
    logic[7:0] _e_1355;
    (* src = "src/generated_driver.spade:364,2" *)
    logic[15:0] _e_1353;
    logic[7:0] _e_1357;
    logic[7:0] _e_1358;
    (* src = "src/generated_driver.spade:365,2" *)
    logic[15:0] _e_1356;
    logic[7:0] _e_1360;
    logic[7:0] _e_1361;
    (* src = "src/generated_driver.spade:366,2" *)
    logic[15:0] _e_1359;
    logic[7:0] _e_1363;
    logic[7:0] _e_1364;
    (* src = "src/generated_driver.spade:367,2" *)
    logic[15:0] _e_1362;
    logic[7:0] _e_1366;
    logic[7:0] _e_1367;
    (* src = "src/generated_driver.spade:368,2" *)
    logic[15:0] _e_1365;
    logic[7:0] _e_1369;
    logic[7:0] _e_1370;
    (* src = "src/generated_driver.spade:369,2" *)
    logic[15:0] _e_1368;
    logic[7:0] _e_1372;
    logic[7:0] _e_1373;
    (* src = "src/generated_driver.spade:370,2" *)
    logic[15:0] _e_1371;
    logic[7:0] _e_1375;
    logic[7:0] _e_1376;
    (* src = "src/generated_driver.spade:371,2" *)
    logic[15:0] _e_1374;
    logic[7:0] _e_1378;
    logic[7:0] _e_1379;
    (* src = "src/generated_driver.spade:372,2" *)
    logic[15:0] _e_1377;
    logic[7:0] _e_1381;
    logic[7:0] _e_1382;
    (* src = "src/generated_driver.spade:373,2" *)
    logic[15:0] _e_1380;
    logic[7:0] _e_1384;
    logic[7:0] _e_1385;
    (* src = "src/generated_driver.spade:374,2" *)
    logic[15:0] _e_1383;
    logic[7:0] _e_1387;
    logic[7:0] _e_1388;
    (* src = "src/generated_driver.spade:375,2" *)
    logic[15:0] _e_1386;
    logic[7:0] _e_1390;
    logic[7:0] _e_1391;
    (* src = "src/generated_driver.spade:376,2" *)
    logic[15:0] _e_1389;
    logic[7:0] _e_1393;
    logic[7:0] _e_1394;
    (* src = "src/generated_driver.spade:377,2" *)
    logic[15:0] _e_1392;
    logic[7:0] _e_1396;
    logic[7:0] _e_1397;
    (* src = "src/generated_driver.spade:378,2" *)
    logic[15:0] _e_1395;
    logic[7:0] _e_1399;
    logic[7:0] _e_1400;
    (* src = "src/generated_driver.spade:379,2" *)
    logic[15:0] _e_1398;
    logic[7:0] _e_1402;
    logic[7:0] _e_1403;
    (* src = "src/generated_driver.spade:380,2" *)
    logic[15:0] _e_1401;
    logic[7:0] _e_1405;
    logic[7:0] _e_1406;
    (* src = "src/generated_driver.spade:381,2" *)
    logic[15:0] _e_1404;
    logic[7:0] _e_1408;
    logic[7:0] _e_1409;
    (* src = "src/generated_driver.spade:382,2" *)
    logic[15:0] _e_1407;
    logic[7:0] _e_1411;
    logic[7:0] _e_1412;
    (* src = "src/generated_driver.spade:383,2" *)
    logic[15:0] _e_1410;
    logic[7:0] _e_1414;
    logic[7:0] _e_1415;
    (* src = "src/generated_driver.spade:384,2" *)
    logic[15:0] _e_1413;
    logic[7:0] _e_1417;
    logic[7:0] _e_1418;
    (* src = "src/generated_driver.spade:385,2" *)
    logic[15:0] _e_1416;
    logic[7:0] _e_1420;
    logic[7:0] _e_1421;
    (* src = "src/generated_driver.spade:386,2" *)
    logic[15:0] _e_1419;
    logic[7:0] _e_1423;
    logic[7:0] _e_1424;
    (* src = "src/generated_driver.spade:387,2" *)
    logic[15:0] _e_1422;
    logic[7:0] _e_1426;
    logic[7:0] _e_1427;
    (* src = "src/generated_driver.spade:388,2" *)
    logic[15:0] _e_1425;
    logic[7:0] _e_1429;
    logic[7:0] _e_1430;
    (* src = "src/generated_driver.spade:389,2" *)
    logic[15:0] _e_1428;
    logic[7:0] _e_1432;
    logic[7:0] _e_1433;
    (* src = "src/generated_driver.spade:390,2" *)
    logic[15:0] _e_1431;
    logic[7:0] _e_1435;
    logic[7:0] _e_1436;
    (* src = "src/generated_driver.spade:391,2" *)
    logic[15:0] _e_1434;
    logic[7:0] _e_1438;
    logic[7:0] _e_1439;
    (* src = "src/generated_driver.spade:392,2" *)
    logic[15:0] _e_1437;
    logic[7:0] _e_1441;
    logic[7:0] _e_1442;
    (* src = "src/generated_driver.spade:393,2" *)
    logic[15:0] _e_1440;
    logic[7:0] _e_1444;
    logic[7:0] _e_1445;
    (* src = "src/generated_driver.spade:394,2" *)
    logic[15:0] _e_1443;
    logic[7:0] _e_1447;
    logic[7:0] _e_1448;
    (* src = "src/generated_driver.spade:395,2" *)
    logic[15:0] _e_1446;
    logic[7:0] _e_1450;
    logic[7:0] _e_1451;
    (* src = "src/generated_driver.spade:396,2" *)
    logic[15:0] _e_1449;
    logic[7:0] _e_1453;
    logic[7:0] _e_1454;
    (* src = "src/generated_driver.spade:397,2" *)
    logic[15:0] _e_1452;
    logic[7:0] _e_1456;
    logic[7:0] _e_1457;
    (* src = "src/generated_driver.spade:398,2" *)
    logic[15:0] _e_1455;
    logic[7:0] _e_1459;
    logic[7:0] _e_1460;
    (* src = "src/generated_driver.spade:399,2" *)
    logic[15:0] _e_1458;
    logic[7:0] _e_1462;
    logic[7:0] _e_1463;
    (* src = "src/generated_driver.spade:400,2" *)
    logic[15:0] _e_1461;
    logic[7:0] _e_1465;
    logic[7:0] _e_1466;
    (* src = "src/generated_driver.spade:401,2" *)
    logic[15:0] _e_1464;
    logic[7:0] _e_1468;
    logic[7:0] _e_1469;
    (* src = "src/generated_driver.spade:402,2" *)
    logic[15:0] _e_1467;
    logic[7:0] _e_1471;
    logic[7:0] _e_1472;
    (* src = "src/generated_driver.spade:403,2" *)
    logic[15:0] _e_1470;
    logic[7:0] _e_1474;
    logic[7:0] _e_1475;
    (* src = "src/generated_driver.spade:404,2" *)
    logic[15:0] _e_1473;
    logic[7:0] _e_1477;
    logic[7:0] _e_1478;
    (* src = "src/generated_driver.spade:405,2" *)
    logic[15:0] _e_1476;
    logic[7:0] _e_1480;
    logic[7:0] _e_1481;
    (* src = "src/generated_driver.spade:406,2" *)
    logic[15:0] _e_1479;
    logic[7:0] _e_1483;
    logic[7:0] _e_1484;
    (* src = "src/generated_driver.spade:407,2" *)
    logic[15:0] _e_1482;
    logic[7:0] _e_1486;
    logic[7:0] _e_1487;
    (* src = "src/generated_driver.spade:408,2" *)
    logic[15:0] _e_1485;
    logic[7:0] _e_1489;
    logic[7:0] _e_1490;
    (* src = "src/generated_driver.spade:409,2" *)
    logic[15:0] _e_1488;
    logic[7:0] _e_1492;
    logic[7:0] _e_1493;
    (* src = "src/generated_driver.spade:410,2" *)
    logic[15:0] _e_1491;
    logic[7:0] _e_1495;
    logic[7:0] _e_1496;
    (* src = "src/generated_driver.spade:411,2" *)
    logic[15:0] _e_1494;
    logic[7:0] _e_1498;
    logic[7:0] _e_1499;
    (* src = "src/generated_driver.spade:412,2" *)
    logic[15:0] _e_1497;
    logic[7:0] _e_1501;
    logic[7:0] _e_1502;
    (* src = "src/generated_driver.spade:413,2" *)
    logic[15:0] _e_1500;
    logic[7:0] _e_1504;
    logic[7:0] _e_1505;
    (* src = "src/generated_driver.spade:414,2" *)
    logic[15:0] _e_1503;
    logic[7:0] _e_1507;
    logic[7:0] _e_1508;
    (* src = "src/generated_driver.spade:415,2" *)
    logic[15:0] _e_1506;
    logic[7:0] _e_1510;
    logic[7:0] _e_1511;
    (* src = "src/generated_driver.spade:416,2" *)
    logic[15:0] _e_1509;
    logic[7:0] _e_1513;
    logic[7:0] _e_1514;
    (* src = "src/generated_driver.spade:417,2" *)
    logic[15:0] _e_1512;
    logic[7:0] _e_1516;
    logic[7:0] _e_1517;
    (* src = "src/generated_driver.spade:418,2" *)
    logic[15:0] _e_1515;
    logic[7:0] _e_1519;
    logic[7:0] _e_1520;
    (* src = "src/generated_driver.spade:419,2" *)
    logic[15:0] _e_1518;
    logic[7:0] _e_1522;
    logic[7:0] _e_1523;
    (* src = "src/generated_driver.spade:420,2" *)
    logic[15:0] _e_1521;
    logic[7:0] _e_1525;
    logic[7:0] _e_1526;
    (* src = "src/generated_driver.spade:421,2" *)
    logic[15:0] _e_1524;
    logic[7:0] _e_1528;
    logic[7:0] _e_1529;
    (* src = "src/generated_driver.spade:422,2" *)
    logic[15:0] _e_1527;
    logic[7:0] _e_1531;
    logic[7:0] _e_1532;
    (* src = "src/generated_driver.spade:423,2" *)
    logic[15:0] _e_1530;
    logic[7:0] _e_1534;
    logic[7:0] _e_1535;
    (* src = "src/generated_driver.spade:424,2" *)
    logic[15:0] _e_1533;
    logic[7:0] _e_1537;
    logic[7:0] _e_1538;
    (* src = "src/generated_driver.spade:425,2" *)
    logic[15:0] _e_1536;
    logic[7:0] _e_1540;
    logic[7:0] _e_1541;
    (* src = "src/generated_driver.spade:426,2" *)
    logic[15:0] _e_1539;
    logic[7:0] _e_1543;
    logic[7:0] _e_1544;
    (* src = "src/generated_driver.spade:427,2" *)
    logic[15:0] _e_1542;
    logic[7:0] _e_1546;
    logic[7:0] _e_1547;
    (* src = "src/generated_driver.spade:428,2" *)
    logic[15:0] _e_1545;
    logic[7:0] _e_1549;
    logic[7:0] _e_1550;
    (* src = "src/generated_driver.spade:429,2" *)
    logic[15:0] _e_1548;
    logic[7:0] _e_1552;
    logic[7:0] _e_1553;
    (* src = "src/generated_driver.spade:430,2" *)
    logic[15:0] _e_1551;
    logic[7:0] _e_1555;
    logic[7:0] _e_1556;
    (* src = "src/generated_driver.spade:431,2" *)
    logic[15:0] _e_1554;
    logic[7:0] _e_1558;
    logic[7:0] _e_1559;
    (* src = "src/generated_driver.spade:432,2" *)
    logic[15:0] _e_1557;
    logic[7:0] _e_1561;
    logic[7:0] _e_1562;
    (* src = "src/generated_driver.spade:433,2" *)
    logic[15:0] _e_1560;
    logic[7:0] _e_1564;
    logic[7:0] _e_1565;
    (* src = "src/generated_driver.spade:434,2" *)
    logic[15:0] _e_1563;
    logic[7:0] _e_1567;
    logic[7:0] _e_1568;
    (* src = "src/generated_driver.spade:435,2" *)
    logic[15:0] _e_1566;
    logic[7:0] _e_1570;
    logic[7:0] _e_1571;
    (* src = "src/generated_driver.spade:436,2" *)
    logic[15:0] _e_1569;
    logic[7:0] _e_1573;
    logic[7:0] _e_1574;
    (* src = "src/generated_driver.spade:437,2" *)
    logic[15:0] _e_1572;
    logic[7:0] _e_1576;
    logic[7:0] _e_1577;
    (* src = "src/generated_driver.spade:438,2" *)
    logic[15:0] _e_1575;
    logic[7:0] _e_1579;
    logic[7:0] _e_1580;
    (* src = "src/generated_driver.spade:439,2" *)
    logic[15:0] _e_1578;
    logic[7:0] _e_1582;
    logic[7:0] _e_1583;
    (* src = "src/generated_driver.spade:440,2" *)
    logic[15:0] _e_1581;
    logic[7:0] _e_1585;
    logic[7:0] _e_1586;
    (* src = "src/generated_driver.spade:441,2" *)
    logic[15:0] _e_1584;
    logic[7:0] _e_1588;
    logic[7:0] _e_1589;
    (* src = "src/generated_driver.spade:442,2" *)
    logic[15:0] _e_1587;
    logic[7:0] _e_1591;
    logic[7:0] _e_1592;
    (* src = "src/generated_driver.spade:443,2" *)
    logic[15:0] _e_1590;
    logic[7:0] _e_1594;
    logic[7:0] _e_1595;
    (* src = "src/generated_driver.spade:444,2" *)
    logic[15:0] _e_1593;
    logic[7:0] _e_1597;
    logic[7:0] _e_1598;
    (* src = "src/generated_driver.spade:445,2" *)
    logic[15:0] _e_1596;
    logic[7:0] _e_1600;
    logic[7:0] _e_1601;
    (* src = "src/generated_driver.spade:446,2" *)
    logic[15:0] _e_1599;
    logic[7:0] _e_1603;
    logic[7:0] _e_1604;
    (* src = "src/generated_driver.spade:447,2" *)
    logic[15:0] _e_1602;
    logic[7:0] _e_1606;
    logic[7:0] _e_1607;
    (* src = "src/generated_driver.spade:448,2" *)
    logic[15:0] _e_1605;
    logic[7:0] _e_1609;
    logic[7:0] _e_1610;
    (* src = "src/generated_driver.spade:449,2" *)
    logic[15:0] _e_1608;
    logic[7:0] _e_1612;
    logic[7:0] _e_1613;
    (* src = "src/generated_driver.spade:450,2" *)
    logic[15:0] _e_1611;
    logic[7:0] _e_1615;
    logic[7:0] _e_1616;
    (* src = "src/generated_driver.spade:451,2" *)
    logic[15:0] _e_1614;
    logic[7:0] _e_1618;
    logic[7:0] _e_1619;
    (* src = "src/generated_driver.spade:452,2" *)
    logic[15:0] _e_1617;
    logic[7:0] _e_1621;
    logic[7:0] _e_1622;
    (* src = "src/generated_driver.spade:453,2" *)
    logic[15:0] _e_1620;
    logic[7:0] _e_1624;
    logic[7:0] _e_1625;
    (* src = "src/generated_driver.spade:454,2" *)
    logic[15:0] _e_1623;
    logic[7:0] _e_1627;
    logic[7:0] _e_1628;
    (* src = "src/generated_driver.spade:455,2" *)
    logic[15:0] _e_1626;
    logic[7:0] _e_1630;
    logic[7:0] _e_1631;
    (* src = "src/generated_driver.spade:456,2" *)
    logic[15:0] _e_1629;
    logic[7:0] _e_1633;
    logic[7:0] _e_1634;
    (* src = "src/generated_driver.spade:457,2" *)
    logic[15:0] _e_1632;
    logic[7:0] _e_1636;
    logic[7:0] _e_1637;
    (* src = "src/generated_driver.spade:458,2" *)
    logic[15:0] _e_1635;
    logic[7:0] _e_1639;
    logic[7:0] _e_1640;
    (* src = "src/generated_driver.spade:459,2" *)
    logic[15:0] _e_1638;
    logic[7:0] _e_1642;
    logic[7:0] _e_1643;
    (* src = "src/generated_driver.spade:460,2" *)
    logic[15:0] _e_1641;
    logic[7:0] _e_1645;
    logic[7:0] _e_1646;
    (* src = "src/generated_driver.spade:461,2" *)
    logic[15:0] _e_1644;
    logic[7:0] _e_1648;
    logic[7:0] _e_1649;
    (* src = "src/generated_driver.spade:462,2" *)
    logic[15:0] _e_1647;
    logic[7:0] _e_1651;
    logic[7:0] _e_1652;
    (* src = "src/generated_driver.spade:463,2" *)
    logic[15:0] _e_1650;
    logic[7:0] _e_1654;
    logic[7:0] _e_1655;
    (* src = "src/generated_driver.spade:464,2" *)
    logic[15:0] _e_1653;
    logic[7:0] _e_1657;
    logic[7:0] _e_1658;
    (* src = "src/generated_driver.spade:465,2" *)
    logic[15:0] _e_1656;
    logic[7:0] _e_1660;
    logic[7:0] _e_1661;
    (* src = "src/generated_driver.spade:466,2" *)
    logic[15:0] _e_1659;
    logic[7:0] _e_1663;
    logic[7:0] _e_1664;
    (* src = "src/generated_driver.spade:467,2" *)
    logic[15:0] _e_1662;
    logic[7:0] _e_1666;
    logic[7:0] _e_1667;
    (* src = "src/generated_driver.spade:468,2" *)
    logic[15:0] _e_1665;
    logic[7:0] _e_1669;
    logic[7:0] _e_1670;
    (* src = "src/generated_driver.spade:469,2" *)
    logic[15:0] _e_1668;
    logic[7:0] _e_1672;
    logic[7:0] _e_1673;
    (* src = "src/generated_driver.spade:470,2" *)
    logic[15:0] _e_1671;
    logic[7:0] _e_1675;
    logic[7:0] _e_1676;
    (* src = "src/generated_driver.spade:471,2" *)
    logic[15:0] _e_1674;
    logic[7:0] _e_1678;
    logic[7:0] _e_1679;
    (* src = "src/generated_driver.spade:472,2" *)
    logic[15:0] _e_1677;
    logic[7:0] _e_1681;
    logic[7:0] _e_1682;
    (* src = "src/generated_driver.spade:473,2" *)
    logic[15:0] _e_1680;
    logic[7:0] _e_1684;
    logic[7:0] _e_1685;
    (* src = "src/generated_driver.spade:474,2" *)
    logic[15:0] _e_1683;
    logic[7:0] _e_1687;
    logic[7:0] _e_1688;
    (* src = "src/generated_driver.spade:475,2" *)
    logic[15:0] _e_1686;
    logic[7:0] _e_1690;
    logic[7:0] _e_1691;
    (* src = "src/generated_driver.spade:476,2" *)
    logic[15:0] _e_1689;
    logic[7:0] _e_1693;
    logic[7:0] _e_1694;
    (* src = "src/generated_driver.spade:477,2" *)
    logic[15:0] _e_1692;
    logic[7:0] _e_1696;
    logic[7:0] _e_1697;
    (* src = "src/generated_driver.spade:478,2" *)
    logic[15:0] _e_1695;
    logic[7:0] _e_1699;
    logic[7:0] _e_1700;
    (* src = "src/generated_driver.spade:479,2" *)
    logic[15:0] _e_1698;
    logic[7:0] _e_1702;
    logic[7:0] _e_1703;
    (* src = "src/generated_driver.spade:480,2" *)
    logic[15:0] _e_1701;
    logic[7:0] _e_1705;
    logic[7:0] _e_1706;
    (* src = "src/generated_driver.spade:481,2" *)
    logic[15:0] _e_1704;
    logic[7:0] _e_1708;
    logic[7:0] _e_1709;
    (* src = "src/generated_driver.spade:482,2" *)
    logic[15:0] _e_1707;
    logic[7:0] _e_1711;
    logic[7:0] _e_1712;
    (* src = "src/generated_driver.spade:483,2" *)
    logic[15:0] _e_1710;
    logic[7:0] _e_1714;
    logic[7:0] _e_1715;
    (* src = "src/generated_driver.spade:484,2" *)
    logic[15:0] _e_1713;
    logic[7:0] _e_1717;
    logic[7:0] _e_1718;
    (* src = "src/generated_driver.spade:485,2" *)
    logic[15:0] _e_1716;
    logic[7:0] _e_1720;
    logic[7:0] _e_1721;
    (* src = "src/generated_driver.spade:486,2" *)
    logic[15:0] _e_1719;
    logic[7:0] _e_1723;
    logic[7:0] _e_1724;
    (* src = "src/generated_driver.spade:487,2" *)
    logic[15:0] _e_1722;
    logic[7:0] _e_1726;
    logic[7:0] _e_1727;
    (* src = "src/generated_driver.spade:488,2" *)
    logic[15:0] _e_1725;
    logic[7:0] _e_1729;
    logic[7:0] _e_1730;
    (* src = "src/generated_driver.spade:489,2" *)
    logic[15:0] _e_1728;
    logic[7:0] _e_1732;
    logic[7:0] _e_1733;
    (* src = "src/generated_driver.spade:490,2" *)
    logic[15:0] _e_1731;
    logic[7:0] _e_1735;
    logic[7:0] _e_1736;
    (* src = "src/generated_driver.spade:491,2" *)
    logic[15:0] _e_1734;
    logic[7:0] _e_1738;
    logic[7:0] _e_1739;
    (* src = "src/generated_driver.spade:492,2" *)
    logic[15:0] _e_1737;
    logic[7:0] _e_1741;
    logic[7:0] _e_1742;
    (* src = "src/generated_driver.spade:493,2" *)
    logic[15:0] _e_1740;
    logic[7:0] _e_1744;
    logic[7:0] _e_1745;
    (* src = "src/generated_driver.spade:494,2" *)
    logic[15:0] _e_1743;
    logic[7:0] _e_1747;
    logic[7:0] _e_1748;
    (* src = "src/generated_driver.spade:495,2" *)
    logic[15:0] _e_1746;
    logic[7:0] _e_1750;
    logic[7:0] _e_1751;
    (* src = "src/generated_driver.spade:496,2" *)
    logic[15:0] _e_1749;
    logic[7:0] _e_1753;
    logic[7:0] _e_1754;
    (* src = "src/generated_driver.spade:497,2" *)
    logic[15:0] _e_1752;
    logic[7:0] _e_1756;
    logic[7:0] _e_1757;
    (* src = "src/generated_driver.spade:498,2" *)
    logic[15:0] _e_1755;
    logic[7:0] _e_1759;
    logic[7:0] _e_1760;
    (* src = "src/generated_driver.spade:499,2" *)
    logic[15:0] _e_1758;
    logic[7:0] _e_1762;
    logic[7:0] _e_1763;
    (* src = "src/generated_driver.spade:500,2" *)
    logic[15:0] _e_1761;
    logic[7:0] _e_1765;
    logic[7:0] _e_1766;
    (* src = "src/generated_driver.spade:501,2" *)
    logic[15:0] _e_1764;
    logic[7:0] _e_1768;
    logic[7:0] _e_1769;
    (* src = "src/generated_driver.spade:502,2" *)
    logic[15:0] _e_1767;
    logic[7:0] _e_1771;
    logic[7:0] _e_1772;
    (* src = "src/generated_driver.spade:503,2" *)
    logic[15:0] _e_1770;
    logic[7:0] _e_1774;
    logic[7:0] _e_1775;
    (* src = "src/generated_driver.spade:504,2" *)
    logic[15:0] _e_1773;
    logic[7:0] _e_1777;
    logic[7:0] _e_1778;
    (* src = "src/generated_driver.spade:505,2" *)
    logic[15:0] _e_1776;
    logic[7:0] _e_1780;
    logic[7:0] _e_1781;
    (* src = "src/generated_driver.spade:506,2" *)
    logic[15:0] _e_1779;
    logic[7:0] _e_1783;
    logic[7:0] _e_1784;
    (* src = "src/generated_driver.spade:507,2" *)
    logic[15:0] _e_1782;
    logic[7:0] _e_1786;
    logic[7:0] _e_1787;
    (* src = "src/generated_driver.spade:508,2" *)
    logic[15:0] _e_1785;
    logic[7:0] _e_1789;
    logic[7:0] _e_1790;
    (* src = "src/generated_driver.spade:509,2" *)
    logic[15:0] _e_1788;
    logic[7:0] _e_1792;
    logic[7:0] _e_1793;
    (* src = "src/generated_driver.spade:510,2" *)
    logic[15:0] _e_1791;
    logic[7:0] _e_1795;
    logic[7:0] _e_1796;
    (* src = "src/generated_driver.spade:511,2" *)
    logic[15:0] _e_1794;
    logic[7:0] _e_1798;
    logic[7:0] _e_1799;
    (* src = "src/generated_driver.spade:512,2" *)
    logic[15:0] _e_1797;
    logic[7:0] _e_1801;
    logic[7:0] _e_1802;
    (* src = "src/generated_driver.spade:513,2" *)
    logic[15:0] _e_1800;
    logic[7:0] _e_1804;
    logic[7:0] _e_1805;
    (* src = "src/generated_driver.spade:514,2" *)
    logic[15:0] _e_1803;
    logic[7:0] _e_1807;
    logic[7:0] _e_1808;
    (* src = "src/generated_driver.spade:515,2" *)
    logic[15:0] _e_1806;
    logic[7:0] _e_1810;
    logic[7:0] _e_1811;
    (* src = "src/generated_driver.spade:516,2" *)
    logic[15:0] _e_1809;
    logic[7:0] _e_1813;
    logic[7:0] _e_1814;
    (* src = "src/generated_driver.spade:517,2" *)
    logic[15:0] _e_1812;
    logic[7:0] _e_1816;
    logic[7:0] _e_1817;
    (* src = "src/generated_driver.spade:518,2" *)
    logic[15:0] _e_1815;
    logic[7:0] _e_1819;
    logic[7:0] _e_1820;
    (* src = "src/generated_driver.spade:519,2" *)
    logic[15:0] _e_1818;
    logic[7:0] _e_1822;
    logic[7:0] _e_1823;
    (* src = "src/generated_driver.spade:520,2" *)
    logic[15:0] _e_1821;
    logic[7:0] _e_1825;
    logic[7:0] _e_1826;
    (* src = "src/generated_driver.spade:521,2" *)
    logic[15:0] _e_1824;
    logic[7:0] _e_1828;
    logic[7:0] _e_1829;
    (* src = "src/generated_driver.spade:522,2" *)
    logic[15:0] _e_1827;
    logic[7:0] _e_1831;
    logic[7:0] _e_1832;
    (* src = "src/generated_driver.spade:523,2" *)
    logic[15:0] _e_1830;
    logic[7:0] _e_1834;
    logic[7:0] _e_1835;
    (* src = "src/generated_driver.spade:524,2" *)
    logic[15:0] _e_1833;
    logic[7:0] _e_1837;
    logic[7:0] _e_1838;
    (* src = "src/generated_driver.spade:525,2" *)
    logic[15:0] _e_1836;
    logic[7:0] _e_1840;
    logic[7:0] _e_1841;
    (* src = "src/generated_driver.spade:526,2" *)
    logic[15:0] _e_1839;
    logic[7:0] _e_1843;
    logic[7:0] _e_1844;
    (* src = "src/generated_driver.spade:527,2" *)
    logic[15:0] _e_1842;
    logic[7:0] _e_1846;
    logic[7:0] _e_1847;
    (* src = "src/generated_driver.spade:528,2" *)
    logic[15:0] _e_1845;
    logic[7:0] _e_1849;
    logic[7:0] _e_1850;
    (* src = "src/generated_driver.spade:529,2" *)
    logic[15:0] _e_1848;
    logic[7:0] _e_1852;
    logic[7:0] _e_1853;
    (* src = "src/generated_driver.spade:530,2" *)
    logic[15:0] _e_1851;
    logic[7:0] _e_1855;
    logic[7:0] _e_1856;
    (* src = "src/generated_driver.spade:531,2" *)
    logic[15:0] _e_1854;
    logic[7:0] _e_1858;
    logic[7:0] _e_1859;
    (* src = "src/generated_driver.spade:532,2" *)
    logic[15:0] _e_1857;
    logic[7:0] _e_1861;
    logic[7:0] _e_1862;
    (* src = "src/generated_driver.spade:533,2" *)
    logic[15:0] _e_1860;
    logic[7:0] _e_1864;
    logic[7:0] _e_1865;
    (* src = "src/generated_driver.spade:534,2" *)
    logic[15:0] _e_1863;
    logic[7:0] _e_1867;
    logic[7:0] _e_1868;
    (* src = "src/generated_driver.spade:535,2" *)
    logic[15:0] _e_1866;
    logic[7:0] _e_1870;
    logic[7:0] _e_1871;
    (* src = "src/generated_driver.spade:536,2" *)
    logic[15:0] _e_1869;
    logic[7:0] _e_1873;
    logic[7:0] _e_1874;
    (* src = "src/generated_driver.spade:537,2" *)
    logic[15:0] _e_1872;
    logic[7:0] _e_1876;
    logic[7:0] _e_1877;
    (* src = "src/generated_driver.spade:538,2" *)
    logic[15:0] _e_1875;
    logic[7:0] _e_1879;
    logic[7:0] _e_1880;
    (* src = "src/generated_driver.spade:539,2" *)
    logic[15:0] _e_1878;
    logic[7:0] _e_1882;
    logic[7:0] _e_1883;
    (* src = "src/generated_driver.spade:540,2" *)
    logic[15:0] _e_1881;
    logic[7:0] _e_1885;
    logic[7:0] _e_1886;
    (* src = "src/generated_driver.spade:541,2" *)
    logic[15:0] _e_1884;
    logic[7:0] _e_1888;
    logic[7:0] _e_1889;
    (* src = "src/generated_driver.spade:542,2" *)
    logic[15:0] _e_1887;
    logic[7:0] _e_1891;
    logic[7:0] _e_1892;
    (* src = "src/generated_driver.spade:543,2" *)
    logic[15:0] _e_1890;
    logic[7:0] _e_1894;
    logic[7:0] _e_1895;
    (* src = "src/generated_driver.spade:544,2" *)
    logic[15:0] _e_1893;
    logic[7:0] _e_1897;
    logic[7:0] _e_1898;
    (* src = "src/generated_driver.spade:545,2" *)
    logic[15:0] _e_1896;
    logic[7:0] _e_1900;
    logic[7:0] _e_1901;
    (* src = "src/generated_driver.spade:546,2" *)
    logic[15:0] _e_1899;
    logic[7:0] _e_1903;
    logic[7:0] _e_1904;
    (* src = "src/generated_driver.spade:547,2" *)
    logic[15:0] _e_1902;
    logic[7:0] _e_1906;
    logic[7:0] _e_1907;
    (* src = "src/generated_driver.spade:548,2" *)
    logic[15:0] _e_1905;
    logic[7:0] _e_1909;
    logic[7:0] _e_1910;
    (* src = "src/generated_driver.spade:549,2" *)
    logic[15:0] _e_1908;
    logic[7:0] _e_1912;
    logic[7:0] _e_1913;
    (* src = "src/generated_driver.spade:550,2" *)
    logic[15:0] _e_1911;
    logic[7:0] _e_1915;
    logic[7:0] _e_1916;
    (* src = "src/generated_driver.spade:551,2" *)
    logic[15:0] _e_1914;
    logic[7:0] _e_1918;
    logic[7:0] _e_1919;
    (* src = "src/generated_driver.spade:552,2" *)
    logic[15:0] _e_1917;
    logic[7:0] _e_1921;
    logic[7:0] _e_1922;
    (* src = "src/generated_driver.spade:553,2" *)
    logic[15:0] _e_1920;
    logic[7:0] _e_1924;
    logic[7:0] _e_1925;
    (* src = "src/generated_driver.spade:554,2" *)
    logic[15:0] _e_1923;
    logic[7:0] _e_1927;
    logic[7:0] _e_1928;
    (* src = "src/generated_driver.spade:555,2" *)
    logic[15:0] _e_1926;
    logic[7:0] _e_1930;
    logic[7:0] _e_1931;
    (* src = "src/generated_driver.spade:556,2" *)
    logic[15:0] _e_1929;
    logic[7:0] _e_1933;
    logic[7:0] _e_1934;
    (* src = "src/generated_driver.spade:557,2" *)
    logic[15:0] _e_1932;
    logic[7:0] _e_1936;
    logic[7:0] _e_1937;
    (* src = "src/generated_driver.spade:558,2" *)
    logic[15:0] _e_1935;
    logic[7:0] _e_1939;
    logic[7:0] _e_1940;
    (* src = "src/generated_driver.spade:559,2" *)
    logic[15:0] _e_1938;
    logic[7:0] _e_1942;
    logic[7:0] _e_1943;
    (* src = "src/generated_driver.spade:560,2" *)
    logic[15:0] _e_1941;
    logic[7:0] _e_1945;
    logic[7:0] _e_1946;
    (* src = "src/generated_driver.spade:561,2" *)
    logic[15:0] _e_1944;
    logic[7:0] _e_1948;
    logic[7:0] _e_1949;
    (* src = "src/generated_driver.spade:562,2" *)
    logic[15:0] _e_1947;
    logic[7:0] _e_1951;
    logic[7:0] _e_1952;
    (* src = "src/generated_driver.spade:563,2" *)
    logic[15:0] _e_1950;
    logic[7:0] _e_1954;
    logic[7:0] _e_1955;
    (* src = "src/generated_driver.spade:564,2" *)
    logic[15:0] _e_1953;
    logic[7:0] _e_1957;
    logic[7:0] _e_1958;
    (* src = "src/generated_driver.spade:565,2" *)
    logic[15:0] _e_1956;
    logic[7:0] _e_1960;
    logic[7:0] _e_1961;
    (* src = "src/generated_driver.spade:566,2" *)
    logic[15:0] _e_1959;
    logic[7:0] _e_1963;
    logic[7:0] _e_1964;
    (* src = "src/generated_driver.spade:567,2" *)
    logic[15:0] _e_1962;
    logic[7:0] _e_1966;
    logic[7:0] _e_1967;
    (* src = "src/generated_driver.spade:568,2" *)
    logic[15:0] _e_1965;
    logic[7:0] _e_1969;
    logic[7:0] _e_1970;
    (* src = "src/generated_driver.spade:569,2" *)
    logic[15:0] _e_1968;
    logic[7:0] _e_1972;
    logic[7:0] _e_1973;
    (* src = "src/generated_driver.spade:570,2" *)
    logic[15:0] _e_1971;
    logic[7:0] _e_1975;
    logic[7:0] _e_1976;
    (* src = "src/generated_driver.spade:571,2" *)
    logic[15:0] _e_1974;
    logic[7:0] _e_1978;
    logic[7:0] _e_1979;
    (* src = "src/generated_driver.spade:572,2" *)
    logic[15:0] _e_1977;
    logic[7:0] _e_1981;
    logic[7:0] _e_1982;
    (* src = "src/generated_driver.spade:573,2" *)
    logic[15:0] _e_1980;
    logic[7:0] _e_1984;
    logic[7:0] _e_1985;
    (* src = "src/generated_driver.spade:574,2" *)
    logic[15:0] _e_1983;
    logic[7:0] _e_1987;
    logic[7:0] _e_1988;
    (* src = "src/generated_driver.spade:575,2" *)
    logic[15:0] _e_1986;
    logic[7:0] _e_1990;
    logic[7:0] _e_1991;
    (* src = "src/generated_driver.spade:576,2" *)
    logic[15:0] _e_1989;
    logic[7:0] _e_1993;
    logic[7:0] _e_1994;
    (* src = "src/generated_driver.spade:577,2" *)
    logic[15:0] _e_1992;
    logic[7:0] _e_1996;
    logic[7:0] _e_1997;
    (* src = "src/generated_driver.spade:578,2" *)
    logic[15:0] _e_1995;
    logic[7:0] _e_1999;
    logic[7:0] _e_2000;
    (* src = "src/generated_driver.spade:579,2" *)
    logic[15:0] _e_1998;
    logic[7:0] _e_2002;
    logic[7:0] _e_2003;
    (* src = "src/generated_driver.spade:580,2" *)
    logic[15:0] _e_2001;
    logic[7:0] _e_2005;
    logic[7:0] _e_2006;
    (* src = "src/generated_driver.spade:581,2" *)
    logic[15:0] _e_2004;
    logic[7:0] _e_2008;
    logic[7:0] _e_2009;
    (* src = "src/generated_driver.spade:582,2" *)
    logic[15:0] _e_2007;
    logic[7:0] _e_2011;
    logic[7:0] _e_2012;
    (* src = "src/generated_driver.spade:583,2" *)
    logic[15:0] _e_2010;
    logic[7:0] _e_2014;
    logic[7:0] _e_2015;
    (* src = "src/generated_driver.spade:584,2" *)
    logic[15:0] _e_2013;
    logic[7:0] _e_2017;
    logic[7:0] _e_2018;
    (* src = "src/generated_driver.spade:585,2" *)
    logic[15:0] _e_2016;
    logic[7:0] _e_2020;
    logic[7:0] _e_2021;
    (* src = "src/generated_driver.spade:586,2" *)
    logic[15:0] _e_2019;
    logic[7:0] _e_2023;
    logic[7:0] _e_2024;
    (* src = "src/generated_driver.spade:587,2" *)
    logic[15:0] _e_2022;
    logic[7:0] _e_2026;
    logic[7:0] _e_2027;
    (* src = "src/generated_driver.spade:588,2" *)
    logic[15:0] _e_2025;
    logic[7:0] _e_2029;
    logic[7:0] _e_2030;
    (* src = "src/generated_driver.spade:589,2" *)
    logic[15:0] _e_2028;
    logic[7:0] _e_2032;
    logic[7:0] _e_2033;
    (* src = "src/generated_driver.spade:590,2" *)
    logic[15:0] _e_2031;
    logic[7:0] _e_2035;
    logic[7:0] _e_2036;
    (* src = "src/generated_driver.spade:591,2" *)
    logic[15:0] _e_2034;
    logic[7:0] _e_2038;
    logic[7:0] _e_2039;
    (* src = "src/generated_driver.spade:592,2" *)
    logic[15:0] _e_2037;
    logic[7:0] _e_2041;
    logic[7:0] _e_2042;
    (* src = "src/generated_driver.spade:593,2" *)
    logic[15:0] _e_2040;
    logic[7:0] _e_2044;
    logic[7:0] _e_2045;
    (* src = "src/generated_driver.spade:594,2" *)
    logic[15:0] _e_2043;
    logic[7:0] _e_2047;
    logic[7:0] _e_2048;
    (* src = "src/generated_driver.spade:595,2" *)
    logic[15:0] _e_2046;
    logic[7:0] _e_2050;
    logic[7:0] _e_2051;
    (* src = "src/generated_driver.spade:596,2" *)
    logic[15:0] _e_2049;
    logic[7:0] _e_2053;
    logic[7:0] _e_2054;
    (* src = "src/generated_driver.spade:597,2" *)
    logic[15:0] _e_2052;
    logic[7:0] _e_2056;
    logic[7:0] _e_2057;
    (* src = "src/generated_driver.spade:598,2" *)
    logic[15:0] _e_2055;
    logic[7:0] _e_2059;
    logic[7:0] _e_2060;
    (* src = "src/generated_driver.spade:599,2" *)
    logic[15:0] _e_2058;
    logic[7:0] _e_2062;
    logic[7:0] _e_2063;
    (* src = "src/generated_driver.spade:600,2" *)
    logic[15:0] _e_2061;
    logic[7:0] _e_2065;
    logic[7:0] _e_2066;
    (* src = "src/generated_driver.spade:601,2" *)
    logic[15:0] _e_2064;
    logic[7:0] _e_2068;
    logic[7:0] _e_2069;
    (* src = "src/generated_driver.spade:602,2" *)
    logic[15:0] _e_2067;
    logic[7:0] _e_2071;
    logic[7:0] _e_2072;
    (* src = "src/generated_driver.spade:603,2" *)
    logic[15:0] _e_2070;
    logic[7:0] _e_2074;
    logic[7:0] _e_2075;
    (* src = "src/generated_driver.spade:604,2" *)
    logic[15:0] _e_2073;
    logic[7:0] _e_2077;
    logic[7:0] _e_2078;
    (* src = "src/generated_driver.spade:605,2" *)
    logic[15:0] _e_2076;
    logic[7:0] _e_2080;
    logic[7:0] _e_2081;
    (* src = "src/generated_driver.spade:606,2" *)
    logic[15:0] _e_2079;
    logic[7:0] _e_2083;
    logic[7:0] _e_2084;
    (* src = "src/generated_driver.spade:607,2" *)
    logic[15:0] _e_2082;
    logic[7:0] _e_2086;
    logic[7:0] _e_2087;
    (* src = "src/generated_driver.spade:608,2" *)
    logic[15:0] _e_2085;
    logic[7:0] _e_2089;
    logic[7:0] _e_2090;
    (* src = "src/generated_driver.spade:609,2" *)
    logic[15:0] _e_2088;
    logic[7:0] _e_2092;
    logic[7:0] _e_2093;
    (* src = "src/generated_driver.spade:610,2" *)
    logic[15:0] _e_2091;
    logic[7:0] _e_2095;
    logic[7:0] _e_2096;
    (* src = "src/generated_driver.spade:611,2" *)
    logic[15:0] _e_2094;
    logic[7:0] _e_2098;
    logic[7:0] _e_2099;
    (* src = "src/generated_driver.spade:612,2" *)
    logic[15:0] _e_2097;
    logic[7:0] _e_2101;
    logic[7:0] _e_2102;
    (* src = "src/generated_driver.spade:613,2" *)
    logic[15:0] _e_2100;
    logic[7:0] _e_2104;
    logic[7:0] _e_2105;
    (* src = "src/generated_driver.spade:614,2" *)
    logic[15:0] _e_2103;
    logic[7:0] _e_2107;
    logic[7:0] _e_2108;
    (* src = "src/generated_driver.spade:615,2" *)
    logic[15:0] _e_2106;
    logic[7:0] _e_2110;
    logic[7:0] _e_2111;
    (* src = "src/generated_driver.spade:616,2" *)
    logic[15:0] _e_2109;
    logic[7:0] _e_2113;
    logic[7:0] _e_2114;
    (* src = "src/generated_driver.spade:617,2" *)
    logic[15:0] _e_2112;
    logic[7:0] _e_2116;
    logic[7:0] _e_2117;
    (* src = "src/generated_driver.spade:618,2" *)
    logic[15:0] _e_2115;
    logic[7:0] _e_2119;
    logic[7:0] _e_2120;
    (* src = "src/generated_driver.spade:619,2" *)
    logic[15:0] _e_2118;
    logic[7:0] _e_2122;
    logic[7:0] _e_2123;
    (* src = "src/generated_driver.spade:620,2" *)
    logic[15:0] _e_2121;
    logic[7:0] _e_2125;
    logic[7:0] _e_2126;
    (* src = "src/generated_driver.spade:621,2" *)
    logic[15:0] _e_2124;
    logic[7:0] _e_2128;
    logic[7:0] _e_2129;
    (* src = "src/generated_driver.spade:622,2" *)
    logic[15:0] _e_2127;
    logic[7:0] _e_2131;
    logic[7:0] _e_2132;
    (* src = "src/generated_driver.spade:623,2" *)
    logic[15:0] _e_2130;
    logic[7:0] _e_2134;
    logic[7:0] _e_2135;
    (* src = "src/generated_driver.spade:624,2" *)
    logic[15:0] _e_2133;
    logic[7:0] _e_2137;
    logic[7:0] _e_2138;
    (* src = "src/generated_driver.spade:625,2" *)
    logic[15:0] _e_2136;
    logic[7:0] _e_2140;
    logic[7:0] _e_2141;
    (* src = "src/generated_driver.spade:626,2" *)
    logic[15:0] _e_2139;
    logic[7:0] _e_2143;
    logic[7:0] _e_2144;
    (* src = "src/generated_driver.spade:627,2" *)
    logic[15:0] _e_2142;
    logic[7:0] _e_2146;
    logic[7:0] _e_2147;
    (* src = "src/generated_driver.spade:628,2" *)
    logic[15:0] _e_2145;
    logic[7:0] _e_2149;
    logic[7:0] _e_2150;
    (* src = "src/generated_driver.spade:629,2" *)
    logic[15:0] _e_2148;
    logic[7:0] _e_2152;
    logic[7:0] _e_2153;
    (* src = "src/generated_driver.spade:630,2" *)
    logic[15:0] _e_2151;
    logic[7:0] _e_2155;
    logic[7:0] _e_2156;
    (* src = "src/generated_driver.spade:631,2" *)
    logic[15:0] _e_2154;
    logic[7:0] _e_2158;
    logic[7:0] _e_2159;
    (* src = "src/generated_driver.spade:632,2" *)
    logic[15:0] _e_2157;
    logic[7:0] _e_2161;
    logic[7:0] _e_2162;
    (* src = "src/generated_driver.spade:633,2" *)
    logic[15:0] _e_2160;
    logic[7:0] _e_2164;
    logic[7:0] _e_2165;
    (* src = "src/generated_driver.spade:634,2" *)
    logic[15:0] _e_2163;
    logic[7:0] _e_2167;
    logic[7:0] _e_2168;
    (* src = "src/generated_driver.spade:635,2" *)
    logic[15:0] _e_2166;
    logic[7:0] _e_2170;
    logic[7:0] _e_2171;
    (* src = "src/generated_driver.spade:636,2" *)
    logic[15:0] _e_2169;
    logic[7:0] _e_2173;
    logic[7:0] _e_2174;
    (* src = "src/generated_driver.spade:637,2" *)
    logic[15:0] _e_2172;
    logic[7:0] _e_2176;
    logic[7:0] _e_2177;
    (* src = "src/generated_driver.spade:638,2" *)
    logic[15:0] _e_2175;
    logic[7:0] _e_2179;
    logic[7:0] _e_2180;
    (* src = "src/generated_driver.spade:639,2" *)
    logic[15:0] _e_2178;
    logic[7:0] _e_2182;
    logic[7:0] _e_2183;
    (* src = "src/generated_driver.spade:640,2" *)
    logic[15:0] _e_2181;
    logic[7:0] _e_2185;
    logic[7:0] _e_2186;
    (* src = "src/generated_driver.spade:641,2" *)
    logic[15:0] _e_2184;
    logic[7:0] _e_2188;
    logic[7:0] _e_2189;
    (* src = "src/generated_driver.spade:642,2" *)
    logic[15:0] _e_2187;
    logic[7:0] _e_2191;
    logic[7:0] _e_2192;
    (* src = "src/generated_driver.spade:643,2" *)
    logic[15:0] _e_2190;
    logic[7:0] _e_2194;
    logic[7:0] _e_2195;
    (* src = "src/generated_driver.spade:644,2" *)
    logic[15:0] _e_2193;
    logic[7:0] _e_2197;
    logic[7:0] _e_2198;
    (* src = "src/generated_driver.spade:645,2" *)
    logic[15:0] _e_2196;
    logic[7:0] _e_2200;
    logic[7:0] _e_2201;
    (* src = "src/generated_driver.spade:646,2" *)
    logic[15:0] _e_2199;
    logic[7:0] _e_2203;
    logic[7:0] _e_2204;
    (* src = "src/generated_driver.spade:647,2" *)
    logic[15:0] _e_2202;
    logic[7:0] _e_2206;
    logic[7:0] _e_2207;
    (* src = "src/generated_driver.spade:648,2" *)
    logic[15:0] _e_2205;
    logic[7:0] _e_2209;
    logic[7:0] _e_2210;
    (* src = "src/generated_driver.spade:649,2" *)
    logic[15:0] _e_2208;
    logic[7:0] _e_2212;
    logic[7:0] _e_2213;
    (* src = "src/generated_driver.spade:650,2" *)
    logic[15:0] _e_2211;
    logic[7:0] _e_2215;
    logic[7:0] _e_2216;
    (* src = "src/generated_driver.spade:651,2" *)
    logic[15:0] _e_2214;
    logic[7:0] _e_2218;
    logic[7:0] _e_2219;
    (* src = "src/generated_driver.spade:652,2" *)
    logic[15:0] _e_2217;
    logic[7:0] _e_2221;
    logic[7:0] _e_2222;
    (* src = "src/generated_driver.spade:653,2" *)
    logic[15:0] _e_2220;
    logic[7:0] _e_2224;
    logic[7:0] _e_2225;
    (* src = "src/generated_driver.spade:654,2" *)
    logic[15:0] _e_2223;
    logic[7:0] _e_2227;
    logic[7:0] _e_2228;
    (* src = "src/generated_driver.spade:655,2" *)
    logic[15:0] _e_2226;
    logic[7:0] _e_2230;
    logic[7:0] _e_2231;
    (* src = "src/generated_driver.spade:656,2" *)
    logic[15:0] _e_2229;
    logic[7:0] _e_2233;
    logic[7:0] _e_2234;
    (* src = "src/generated_driver.spade:657,2" *)
    logic[15:0] _e_2232;
    logic[7:0] _e_2236;
    logic[7:0] _e_2237;
    (* src = "src/generated_driver.spade:658,2" *)
    logic[15:0] _e_2235;
    logic[7:0] _e_2239;
    logic[7:0] _e_2240;
    (* src = "src/generated_driver.spade:659,2" *)
    logic[15:0] _e_2238;
    logic[7:0] _e_2242;
    logic[7:0] _e_2243;
    (* src = "src/generated_driver.spade:660,2" *)
    logic[15:0] _e_2241;
    logic[7:0] _e_2245;
    logic[7:0] _e_2246;
    (* src = "src/generated_driver.spade:661,2" *)
    logic[15:0] _e_2244;
    logic[7:0] _e_2248;
    logic[7:0] _e_2249;
    (* src = "src/generated_driver.spade:662,2" *)
    logic[15:0] _e_2247;
    logic[7:0] _e_2251;
    logic[7:0] _e_2252;
    (* src = "src/generated_driver.spade:663,2" *)
    logic[15:0] _e_2250;
    logic[7:0] _e_2254;
    logic[7:0] _e_2255;
    (* src = "src/generated_driver.spade:664,2" *)
    logic[15:0] _e_2253;
    logic[7:0] _e_2257;
    logic[7:0] _e_2258;
    (* src = "src/generated_driver.spade:665,2" *)
    logic[15:0] _e_2256;
    logic[7:0] _e_2260;
    logic[7:0] _e_2261;
    (* src = "src/generated_driver.spade:666,2" *)
    logic[15:0] _e_2259;
    logic[7:0] _e_2263;
    logic[7:0] _e_2264;
    (* src = "src/generated_driver.spade:667,2" *)
    logic[15:0] _e_2262;
    logic[7:0] _e_2266;
    logic[7:0] _e_2267;
    (* src = "src/generated_driver.spade:668,2" *)
    logic[15:0] _e_2265;
    logic[7:0] _e_2269;
    logic[7:0] _e_2270;
    (* src = "src/generated_driver.spade:669,2" *)
    logic[15:0] _e_2268;
    logic[7:0] _e_2272;
    logic[7:0] _e_2273;
    (* src = "src/generated_driver.spade:670,2" *)
    logic[15:0] _e_2271;
    logic[7:0] _e_2275;
    logic[7:0] _e_2276;
    (* src = "src/generated_driver.spade:671,2" *)
    logic[15:0] _e_2274;
    logic[7:0] _e_2278;
    logic[7:0] _e_2279;
    (* src = "src/generated_driver.spade:672,2" *)
    logic[15:0] _e_2277;
    logic[7:0] _e_2281;
    logic[7:0] _e_2282;
    (* src = "src/generated_driver.spade:673,2" *)
    logic[15:0] _e_2280;
    logic[7:0] _e_2284;
    logic[7:0] _e_2285;
    (* src = "src/generated_driver.spade:674,2" *)
    logic[15:0] _e_2283;
    logic[7:0] _e_2287;
    logic[7:0] _e_2288;
    (* src = "src/generated_driver.spade:675,2" *)
    logic[15:0] _e_2286;
    logic[7:0] _e_2290;
    logic[7:0] _e_2291;
    (* src = "src/generated_driver.spade:676,2" *)
    logic[15:0] _e_2289;
    logic[7:0] _e_2293;
    logic[7:0] _e_2294;
    (* src = "src/generated_driver.spade:677,2" *)
    logic[15:0] _e_2292;
    logic[7:0] _e_2296;
    logic[7:0] _e_2297;
    (* src = "src/generated_driver.spade:678,2" *)
    logic[15:0] _e_2295;
    logic[7:0] _e_2299;
    logic[7:0] _e_2300;
    (* src = "src/generated_driver.spade:679,2" *)
    logic[15:0] _e_2298;
    logic[7:0] _e_2302;
    logic[7:0] _e_2303;
    (* src = "src/generated_driver.spade:680,2" *)
    logic[15:0] _e_2301;
    logic[7:0] _e_2305;
    logic[7:0] _e_2306;
    (* src = "src/generated_driver.spade:681,2" *)
    logic[15:0] _e_2304;
    logic[7:0] _e_2308;
    logic[7:0] _e_2309;
    (* src = "src/generated_driver.spade:682,2" *)
    logic[15:0] _e_2307;
    logic[7:0] _e_2311;
    logic[7:0] _e_2312;
    (* src = "src/generated_driver.spade:683,2" *)
    logic[15:0] _e_2310;
    logic[7:0] _e_2314;
    logic[7:0] _e_2315;
    (* src = "src/generated_driver.spade:684,2" *)
    logic[15:0] _e_2313;
    logic[7:0] _e_2317;
    logic[7:0] _e_2318;
    (* src = "src/generated_driver.spade:685,2" *)
    logic[15:0] _e_2316;
    logic[7:0] _e_2320;
    logic[7:0] _e_2321;
    (* src = "src/generated_driver.spade:686,2" *)
    logic[15:0] _e_2319;
    logic[7:0] _e_2323;
    logic[7:0] _e_2324;
    (* src = "src/generated_driver.spade:687,2" *)
    logic[15:0] _e_2322;
    logic[7:0] _e_2326;
    logic[7:0] _e_2327;
    (* src = "src/generated_driver.spade:688,2" *)
    logic[15:0] _e_2325;
    logic[7:0] _e_2329;
    logic[7:0] _e_2330;
    (* src = "src/generated_driver.spade:689,2" *)
    logic[15:0] _e_2328;
    logic[7:0] _e_2332;
    logic[7:0] _e_2333;
    (* src = "src/generated_driver.spade:690,2" *)
    logic[15:0] _e_2331;
    logic[7:0] _e_2335;
    logic[7:0] _e_2336;
    (* src = "src/generated_driver.spade:691,2" *)
    logic[15:0] _e_2334;
    logic[7:0] _e_2338;
    logic[7:0] _e_2339;
    (* src = "src/generated_driver.spade:692,2" *)
    logic[15:0] _e_2337;
    logic[7:0] _e_2341;
    logic[7:0] _e_2342;
    (* src = "src/generated_driver.spade:693,2" *)
    logic[15:0] _e_2340;
    logic[7:0] _e_2344;
    logic[7:0] _e_2345;
    (* src = "src/generated_driver.spade:694,2" *)
    logic[15:0] _e_2343;
    logic[7:0] _e_2347;
    logic[7:0] _e_2348;
    (* src = "src/generated_driver.spade:695,2" *)
    logic[15:0] _e_2346;
    logic[7:0] _e_2350;
    logic[7:0] _e_2351;
    (* src = "src/generated_driver.spade:696,2" *)
    logic[15:0] _e_2349;
    logic[7:0] _e_2353;
    logic[7:0] _e_2354;
    (* src = "src/generated_driver.spade:697,2" *)
    logic[15:0] _e_2352;
    logic[7:0] _e_2356;
    logic[7:0] _e_2357;
    (* src = "src/generated_driver.spade:698,2" *)
    logic[15:0] _e_2355;
    logic[7:0] _e_2359;
    logic[7:0] _e_2360;
    (* src = "src/generated_driver.spade:699,2" *)
    logic[15:0] _e_2358;
    logic[7:0] _e_2362;
    logic[7:0] _e_2363;
    (* src = "src/generated_driver.spade:700,2" *)
    logic[15:0] _e_2361;
    logic[7:0] _e_2365;
    logic[7:0] _e_2366;
    (* src = "src/generated_driver.spade:701,2" *)
    logic[15:0] _e_2364;
    logic[7:0] _e_2368;
    logic[7:0] _e_2369;
    (* src = "src/generated_driver.spade:702,2" *)
    logic[15:0] _e_2367;
    logic[7:0] _e_2371;
    logic[7:0] _e_2372;
    (* src = "src/generated_driver.spade:703,2" *)
    logic[15:0] _e_2370;
    logic[7:0] _e_2374;
    logic[7:0] _e_2375;
    (* src = "src/generated_driver.spade:704,2" *)
    logic[15:0] _e_2373;
    logic[7:0] _e_2377;
    logic[7:0] _e_2378;
    (* src = "src/generated_driver.spade:705,2" *)
    logic[15:0] _e_2376;
    logic[7:0] _e_2380;
    logic[7:0] _e_2381;
    (* src = "src/generated_driver.spade:706,2" *)
    logic[15:0] _e_2379;
    logic[7:0] _e_2383;
    logic[7:0] _e_2384;
    (* src = "src/generated_driver.spade:707,2" *)
    logic[15:0] _e_2382;
    logic[7:0] _e_2386;
    logic[7:0] _e_2387;
    (* src = "src/generated_driver.spade:708,2" *)
    logic[15:0] _e_2385;
    logic[7:0] _e_2389;
    logic[7:0] _e_2390;
    (* src = "src/generated_driver.spade:709,2" *)
    logic[15:0] _e_2388;
    logic[7:0] _e_2392;
    logic[7:0] _e_2393;
    (* src = "src/generated_driver.spade:710,2" *)
    logic[15:0] _e_2391;
    logic[7:0] _e_2395;
    logic[7:0] _e_2396;
    (* src = "src/generated_driver.spade:711,2" *)
    logic[15:0] _e_2394;
    logic[7:0] _e_2398;
    logic[7:0] _e_2399;
    (* src = "src/generated_driver.spade:712,2" *)
    logic[15:0] _e_2397;
    logic[7:0] _e_2401;
    logic[7:0] _e_2402;
    (* src = "src/generated_driver.spade:713,2" *)
    logic[15:0] _e_2400;
    logic[7:0] _e_2404;
    logic[7:0] _e_2405;
    (* src = "src/generated_driver.spade:714,2" *)
    logic[15:0] _e_2403;
    logic[7:0] _e_2407;
    logic[7:0] _e_2408;
    (* src = "src/generated_driver.spade:715,2" *)
    logic[15:0] _e_2406;
    logic[7:0] _e_2410;
    logic[7:0] _e_2411;
    (* src = "src/generated_driver.spade:716,2" *)
    logic[15:0] _e_2409;
    logic[7:0] _e_2413;
    logic[7:0] _e_2414;
    (* src = "src/generated_driver.spade:717,2" *)
    logic[15:0] _e_2412;
    logic[7:0] _e_2416;
    logic[7:0] _e_2417;
    (* src = "src/generated_driver.spade:718,2" *)
    logic[15:0] _e_2415;
    logic[7:0] _e_2419;
    logic[7:0] _e_2420;
    (* src = "src/generated_driver.spade:719,2" *)
    logic[15:0] _e_2418;
    logic[7:0] _e_2422;
    logic[7:0] _e_2423;
    (* src = "src/generated_driver.spade:720,2" *)
    logic[15:0] _e_2421;
    logic[7:0] _e_2425;
    logic[7:0] _e_2426;
    (* src = "src/generated_driver.spade:721,2" *)
    logic[15:0] _e_2424;
    logic[7:0] _e_2428;
    logic[7:0] _e_2429;
    (* src = "src/generated_driver.spade:722,2" *)
    logic[15:0] _e_2427;
    logic[7:0] _e_2431;
    logic[7:0] _e_2432;
    (* src = "src/generated_driver.spade:723,2" *)
    logic[15:0] _e_2430;
    logic[7:0] _e_2434;
    logic[7:0] _e_2435;
    (* src = "src/generated_driver.spade:724,2" *)
    logic[15:0] _e_2433;
    logic[7:0] _e_2437;
    logic[7:0] _e_2438;
    (* src = "src/generated_driver.spade:725,2" *)
    logic[15:0] _e_2436;
    logic[7:0] _e_2440;
    logic[7:0] _e_2441;
    (* src = "src/generated_driver.spade:726,2" *)
    logic[15:0] _e_2439;
    logic[7:0] _e_2443;
    logic[7:0] _e_2444;
    (* src = "src/generated_driver.spade:727,2" *)
    logic[15:0] _e_2442;
    logic[7:0] _e_2446;
    logic[7:0] _e_2447;
    (* src = "src/generated_driver.spade:728,2" *)
    logic[15:0] _e_2445;
    logic[7:0] _e_2449;
    logic[7:0] _e_2450;
    (* src = "src/generated_driver.spade:729,2" *)
    logic[15:0] _e_2448;
    logic[7:0] _e_2452;
    logic[7:0] _e_2453;
    (* src = "src/generated_driver.spade:730,2" *)
    logic[15:0] _e_2451;
    logic[7:0] _e_2455;
    logic[7:0] _e_2456;
    (* src = "src/generated_driver.spade:731,2" *)
    logic[15:0] _e_2454;
    logic[7:0] _e_2458;
    logic[7:0] _e_2459;
    (* src = "src/generated_driver.spade:732,2" *)
    logic[15:0] _e_2457;
    logic[7:0] _e_2461;
    logic[7:0] _e_2462;
    (* src = "src/generated_driver.spade:733,2" *)
    logic[15:0] _e_2460;
    logic[7:0] _e_2464;
    logic[7:0] _e_2465;
    (* src = "src/generated_driver.spade:734,2" *)
    logic[15:0] _e_2463;
    logic[7:0] _e_2467;
    logic[7:0] _e_2468;
    (* src = "src/generated_driver.spade:735,2" *)
    logic[15:0] _e_2466;
    logic[7:0] _e_2470;
    logic[7:0] _e_2471;
    (* src = "src/generated_driver.spade:736,2" *)
    logic[15:0] _e_2469;
    logic[7:0] _e_2473;
    logic[7:0] _e_2474;
    (* src = "src/generated_driver.spade:737,2" *)
    logic[15:0] _e_2472;
    logic[7:0] _e_2476;
    logic[7:0] _e_2477;
    (* src = "src/generated_driver.spade:738,2" *)
    logic[15:0] _e_2475;
    logic[7:0] _e_2479;
    logic[7:0] _e_2480;
    (* src = "src/generated_driver.spade:739,2" *)
    logic[15:0] _e_2478;
    logic[7:0] _e_2482;
    logic[7:0] _e_2483;
    (* src = "src/generated_driver.spade:740,2" *)
    logic[15:0] _e_2481;
    logic[7:0] _e_2485;
    logic[7:0] _e_2486;
    (* src = "src/generated_driver.spade:741,2" *)
    logic[15:0] _e_2484;
    logic[7:0] _e_2488;
    logic[7:0] _e_2489;
    (* src = "src/generated_driver.spade:742,2" *)
    logic[15:0] _e_2487;
    logic[7:0] _e_2491;
    logic[7:0] _e_2492;
    (* src = "src/generated_driver.spade:743,2" *)
    logic[15:0] _e_2490;
    logic[7:0] _e_2494;
    logic[7:0] _e_2495;
    (* src = "src/generated_driver.spade:744,2" *)
    logic[15:0] _e_2493;
    logic[7:0] _e_2497;
    logic[7:0] _e_2498;
    (* src = "src/generated_driver.spade:745,2" *)
    logic[15:0] _e_2496;
    logic[7:0] _e_2500;
    logic[7:0] _e_2501;
    (* src = "src/generated_driver.spade:746,2" *)
    logic[15:0] _e_2499;
    logic[7:0] _e_2503;
    logic[7:0] _e_2504;
    (* src = "src/generated_driver.spade:747,2" *)
    logic[15:0] _e_2502;
    logic[7:0] _e_2506;
    logic[7:0] _e_2507;
    (* src = "src/generated_driver.spade:748,2" *)
    logic[15:0] _e_2505;
    logic[7:0] _e_2509;
    logic[7:0] _e_2510;
    (* src = "src/generated_driver.spade:749,2" *)
    logic[15:0] _e_2508;
    logic[7:0] _e_2512;
    logic[7:0] _e_2513;
    (* src = "src/generated_driver.spade:750,2" *)
    logic[15:0] _e_2511;
    logic[7:0] _e_2515;
    logic[7:0] _e_2516;
    (* src = "src/generated_driver.spade:751,2" *)
    logic[15:0] _e_2514;
    logic[7:0] _e_2518;
    logic[7:0] _e_2519;
    (* src = "src/generated_driver.spade:752,2" *)
    logic[15:0] _e_2517;
    logic[7:0] _e_2521;
    logic[7:0] _e_2522;
    (* src = "src/generated_driver.spade:753,2" *)
    logic[15:0] _e_2520;
    logic[7:0] _e_2524;
    logic[7:0] _e_2525;
    (* src = "src/generated_driver.spade:754,2" *)
    logic[15:0] _e_2523;
    logic[7:0] _e_2527;
    logic[7:0] _e_2528;
    (* src = "src/generated_driver.spade:755,2" *)
    logic[15:0] _e_2526;
    logic[7:0] _e_2530;
    logic[7:0] _e_2531;
    (* src = "src/generated_driver.spade:756,2" *)
    logic[15:0] _e_2529;
    logic[7:0] _e_2533;
    logic[7:0] _e_2534;
    (* src = "src/generated_driver.spade:757,2" *)
    logic[15:0] _e_2532;
    logic[7:0] _e_2536;
    logic[7:0] _e_2537;
    (* src = "src/generated_driver.spade:758,2" *)
    logic[15:0] _e_2535;
    logic[7:0] _e_2539;
    logic[7:0] _e_2540;
    (* src = "src/generated_driver.spade:759,2" *)
    logic[15:0] _e_2538;
    logic[7:0] _e_2542;
    logic[7:0] _e_2543;
    (* src = "src/generated_driver.spade:760,2" *)
    logic[15:0] _e_2541;
    logic[7:0] _e_2545;
    logic[7:0] _e_2546;
    (* src = "src/generated_driver.spade:761,2" *)
    logic[15:0] _e_2544;
    logic[7:0] _e_2548;
    logic[7:0] _e_2549;
    (* src = "src/generated_driver.spade:762,2" *)
    logic[15:0] _e_2547;
    logic[7:0] _e_2551;
    logic[7:0] _e_2552;
    (* src = "src/generated_driver.spade:763,2" *)
    logic[15:0] _e_2550;
    logic[7:0] _e_2554;
    logic[7:0] _e_2555;
    (* src = "src/generated_driver.spade:764,2" *)
    logic[15:0] _e_2553;
    logic[7:0] _e_2557;
    logic[7:0] _e_2558;
    (* src = "src/generated_driver.spade:765,2" *)
    logic[15:0] _e_2556;
    logic[7:0] _e_2560;
    logic[7:0] _e_2561;
    (* src = "src/generated_driver.spade:766,2" *)
    logic[15:0] _e_2559;
    logic[7:0] _e_2563;
    logic[7:0] _e_2564;
    (* src = "src/generated_driver.spade:767,2" *)
    logic[15:0] _e_2562;
    logic[7:0] _e_2566;
    logic[7:0] _e_2567;
    (* src = "src/generated_driver.spade:768,2" *)
    logic[15:0] _e_2565;
    logic[7:0] _e_2569;
    logic[7:0] _e_2570;
    (* src = "src/generated_driver.spade:769,2" *)
    logic[15:0] _e_2568;
    logic[7:0] _e_2572;
    logic[7:0] _e_2573;
    (* src = "src/generated_driver.spade:770,2" *)
    logic[15:0] _e_2571;
    logic[7:0] _e_2575;
    logic[7:0] _e_2576;
    (* src = "src/generated_driver.spade:771,2" *)
    logic[15:0] _e_2574;
    logic[7:0] _e_2578;
    logic[7:0] _e_2579;
    (* src = "src/generated_driver.spade:772,2" *)
    logic[15:0] _e_2577;
    logic[7:0] _e_2581;
    logic[7:0] _e_2582;
    (* src = "src/generated_driver.spade:773,2" *)
    logic[15:0] _e_2580;
    logic[7:0] _e_2584;
    logic[7:0] _e_2585;
    (* src = "src/generated_driver.spade:774,2" *)
    logic[15:0] _e_2583;
    logic[7:0] _e_2587;
    logic[7:0] _e_2588;
    (* src = "src/generated_driver.spade:775,2" *)
    logic[15:0] _e_2586;
    logic[7:0] _e_2590;
    logic[7:0] _e_2591;
    (* src = "src/generated_driver.spade:776,2" *)
    logic[15:0] _e_2589;
    logic[7:0] _e_2593;
    logic[7:0] _e_2594;
    (* src = "src/generated_driver.spade:777,2" *)
    logic[15:0] _e_2592;
    logic[7:0] _e_2596;
    logic[7:0] _e_2597;
    (* src = "src/generated_driver.spade:778,2" *)
    logic[15:0] _e_2595;
    logic[7:0] _e_2599;
    logic[7:0] _e_2600;
    (* src = "src/generated_driver.spade:779,2" *)
    logic[15:0] _e_2598;
    logic[7:0] _e_2602;
    logic[7:0] _e_2603;
    (* src = "src/generated_driver.spade:780,2" *)
    logic[15:0] _e_2601;
    logic[7:0] _e_2605;
    logic[7:0] _e_2606;
    (* src = "src/generated_driver.spade:781,2" *)
    logic[15:0] _e_2604;
    logic[7:0] _e_2608;
    logic[7:0] _e_2609;
    (* src = "src/generated_driver.spade:782,2" *)
    logic[15:0] _e_2607;
    logic[7:0] _e_2611;
    logic[7:0] _e_2612;
    (* src = "src/generated_driver.spade:783,2" *)
    logic[15:0] _e_2610;
    logic[7:0] _e_2614;
    logic[7:0] _e_2615;
    (* src = "src/generated_driver.spade:784,2" *)
    logic[15:0] _e_2613;
    logic[7:0] _e_2617;
    logic[7:0] _e_2618;
    (* src = "src/generated_driver.spade:785,2" *)
    logic[15:0] _e_2616;
    logic[7:0] _e_2620;
    logic[7:0] _e_2621;
    (* src = "src/generated_driver.spade:786,2" *)
    logic[15:0] _e_2619;
    logic[7:0] _e_2623;
    logic[7:0] _e_2624;
    (* src = "src/generated_driver.spade:787,2" *)
    logic[15:0] _e_2622;
    logic[7:0] _e_2626;
    logic[7:0] _e_2627;
    (* src = "src/generated_driver.spade:788,2" *)
    logic[15:0] _e_2625;
    logic[7:0] _e_2629;
    logic[7:0] _e_2630;
    (* src = "src/generated_driver.spade:789,2" *)
    logic[15:0] _e_2628;
    logic[7:0] _e_2632;
    logic[7:0] _e_2633;
    (* src = "src/generated_driver.spade:790,2" *)
    logic[15:0] _e_2631;
    logic[7:0] _e_2635;
    logic[7:0] _e_2636;
    (* src = "src/generated_driver.spade:791,2" *)
    logic[15:0] _e_2634;
    logic[7:0] _e_2638;
    logic[7:0] _e_2639;
    (* src = "src/generated_driver.spade:792,2" *)
    logic[15:0] _e_2637;
    logic[7:0] _e_2641;
    logic[7:0] _e_2642;
    (* src = "src/generated_driver.spade:793,2" *)
    logic[15:0] _e_2640;
    logic[7:0] _e_2644;
    logic[7:0] _e_2645;
    (* src = "src/generated_driver.spade:794,2" *)
    logic[15:0] _e_2643;
    logic[7:0] _e_2647;
    logic[7:0] _e_2648;
    (* src = "src/generated_driver.spade:795,2" *)
    logic[15:0] _e_2646;
    logic[7:0] _e_2650;
    logic[7:0] _e_2651;
    (* src = "src/generated_driver.spade:796,2" *)
    logic[15:0] _e_2649;
    logic[7:0] _e_2653;
    logic[7:0] _e_2654;
    (* src = "src/generated_driver.spade:797,2" *)
    logic[15:0] _e_2652;
    logic[7:0] _e_2656;
    logic[7:0] _e_2657;
    (* src = "src/generated_driver.spade:798,2" *)
    logic[15:0] _e_2655;
    logic[7:0] _e_2659;
    logic[7:0] _e_2660;
    (* src = "src/generated_driver.spade:799,2" *)
    logic[15:0] _e_2658;
    logic[7:0] _e_2662;
    logic[7:0] _e_2663;
    (* src = "src/generated_driver.spade:800,2" *)
    logic[15:0] _e_2661;
    logic[7:0] _e_2665;
    logic[7:0] _e_2666;
    (* src = "src/generated_driver.spade:801,2" *)
    logic[15:0] _e_2664;
    logic[7:0] _e_2668;
    logic[7:0] _e_2669;
    (* src = "src/generated_driver.spade:802,2" *)
    logic[15:0] _e_2667;
    logic[7:0] _e_2671;
    logic[7:0] _e_2672;
    (* src = "src/generated_driver.spade:803,2" *)
    logic[15:0] _e_2670;
    logic[7:0] _e_2674;
    logic[7:0] _e_2675;
    (* src = "src/generated_driver.spade:804,2" *)
    logic[15:0] _e_2673;
    logic[7:0] _e_2677;
    logic[7:0] _e_2678;
    (* src = "src/generated_driver.spade:805,2" *)
    logic[15:0] _e_2676;
    logic[7:0] _e_2680;
    logic[7:0] _e_2681;
    (* src = "src/generated_driver.spade:806,2" *)
    logic[15:0] _e_2679;
    logic[7:0] _e_2683;
    logic[7:0] _e_2684;
    (* src = "src/generated_driver.spade:807,2" *)
    logic[15:0] _e_2682;
    logic[7:0] _e_2686;
    logic[7:0] _e_2687;
    (* src = "src/generated_driver.spade:808,2" *)
    logic[15:0] _e_2685;
    logic[7:0] _e_2689;
    logic[7:0] _e_2690;
    (* src = "src/generated_driver.spade:809,2" *)
    logic[15:0] _e_2688;
    logic[7:0] _e_2692;
    logic[7:0] _e_2693;
    (* src = "src/generated_driver.spade:810,2" *)
    logic[15:0] _e_2691;
    logic[7:0] _e_2695;
    logic[7:0] _e_2696;
    (* src = "src/generated_driver.spade:811,2" *)
    logic[15:0] _e_2694;
    logic[7:0] _e_2698;
    logic[7:0] _e_2699;
    (* src = "src/generated_driver.spade:812,2" *)
    logic[15:0] _e_2697;
    logic[7:0] _e_2701;
    logic[7:0] _e_2702;
    (* src = "src/generated_driver.spade:813,2" *)
    logic[15:0] _e_2700;
    logic[7:0] _e_2704;
    logic[7:0] _e_2705;
    (* src = "src/generated_driver.spade:814,2" *)
    logic[15:0] _e_2703;
    logic[7:0] _e_2707;
    logic[7:0] _e_2708;
    (* src = "src/generated_driver.spade:815,2" *)
    logic[15:0] _e_2706;
    logic[7:0] _e_2710;
    logic[7:0] _e_2711;
    (* src = "src/generated_driver.spade:816,2" *)
    logic[15:0] _e_2709;
    logic[7:0] _e_2713;
    logic[7:0] _e_2714;
    (* src = "src/generated_driver.spade:817,2" *)
    logic[15:0] _e_2712;
    logic[7:0] _e_2716;
    logic[7:0] _e_2717;
    (* src = "src/generated_driver.spade:818,2" *)
    logic[15:0] _e_2715;
    logic[7:0] _e_2719;
    logic[7:0] _e_2720;
    (* src = "src/generated_driver.spade:819,2" *)
    logic[15:0] _e_2718;
    logic[7:0] _e_2722;
    logic[7:0] _e_2723;
    (* src = "src/generated_driver.spade:820,2" *)
    logic[15:0] _e_2721;
    logic[7:0] _e_2725;
    logic[7:0] _e_2726;
    (* src = "src/generated_driver.spade:821,2" *)
    logic[15:0] _e_2724;
    logic[7:0] _e_2728;
    logic[7:0] _e_2729;
    (* src = "src/generated_driver.spade:822,2" *)
    logic[15:0] _e_2727;
    logic[7:0] _e_2731;
    logic[7:0] _e_2732;
    (* src = "src/generated_driver.spade:823,2" *)
    logic[15:0] _e_2730;
    logic[7:0] _e_2734;
    logic[7:0] _e_2735;
    (* src = "src/generated_driver.spade:824,2" *)
    logic[15:0] _e_2733;
    logic[7:0] _e_2737;
    logic[7:0] _e_2738;
    (* src = "src/generated_driver.spade:825,2" *)
    logic[15:0] _e_2736;
    logic[7:0] _e_2740;
    logic[7:0] _e_2741;
    (* src = "src/generated_driver.spade:826,2" *)
    logic[15:0] _e_2739;
    logic[7:0] _e_2743;
    logic[7:0] _e_2744;
    (* src = "src/generated_driver.spade:827,2" *)
    logic[15:0] _e_2742;
    logic[7:0] _e_2746;
    logic[7:0] _e_2747;
    (* src = "src/generated_driver.spade:828,2" *)
    logic[15:0] _e_2745;
    logic[7:0] _e_2749;
    logic[7:0] _e_2750;
    (* src = "src/generated_driver.spade:829,2" *)
    logic[15:0] _e_2748;
    logic[7:0] _e_2752;
    logic[7:0] _e_2753;
    (* src = "src/generated_driver.spade:830,2" *)
    logic[15:0] _e_2751;
    logic[7:0] _e_2755;
    logic[7:0] _e_2756;
    (* src = "src/generated_driver.spade:831,2" *)
    logic[15:0] _e_2754;
    logic[7:0] _e_2758;
    logic[7:0] _e_2759;
    (* src = "src/generated_driver.spade:832,2" *)
    logic[15:0] _e_2757;
    logic[7:0] _e_2761;
    logic[7:0] _e_2762;
    (* src = "src/generated_driver.spade:833,2" *)
    logic[15:0] _e_2760;
    logic[7:0] _e_2764;
    logic[7:0] _e_2765;
    (* src = "src/generated_driver.spade:834,2" *)
    logic[15:0] _e_2763;
    logic[7:0] _e_2767;
    logic[7:0] _e_2768;
    (* src = "src/generated_driver.spade:835,2" *)
    logic[15:0] _e_2766;
    logic[7:0] _e_2770;
    logic[7:0] _e_2771;
    (* src = "src/generated_driver.spade:836,2" *)
    logic[15:0] _e_2769;
    logic[7:0] _e_2773;
    logic[7:0] _e_2774;
    (* src = "src/generated_driver.spade:837,2" *)
    logic[15:0] _e_2772;
    logic[7:0] _e_2776;
    logic[7:0] _e_2777;
    (* src = "src/generated_driver.spade:838,2" *)
    logic[15:0] _e_2775;
    logic[7:0] _e_2779;
    logic[7:0] _e_2780;
    (* src = "src/generated_driver.spade:839,2" *)
    logic[15:0] _e_2778;
    logic[7:0] _e_2782;
    logic[7:0] _e_2783;
    (* src = "src/generated_driver.spade:840,2" *)
    logic[15:0] _e_2781;
    logic[7:0] _e_2785;
    logic[7:0] _e_2786;
    (* src = "src/generated_driver.spade:841,2" *)
    logic[15:0] _e_2784;
    logic[7:0] _e_2788;
    logic[7:0] _e_2789;
    (* src = "src/generated_driver.spade:842,2" *)
    logic[15:0] _e_2787;
    logic[7:0] _e_2791;
    logic[7:0] _e_2792;
    (* src = "src/generated_driver.spade:843,2" *)
    logic[15:0] _e_2790;
    logic[7:0] _e_2794;
    logic[7:0] _e_2795;
    (* src = "src/generated_driver.spade:844,2" *)
    logic[15:0] _e_2793;
    logic[7:0] _e_2797;
    logic[7:0] _e_2798;
    (* src = "src/generated_driver.spade:845,2" *)
    logic[15:0] _e_2796;
    logic[7:0] _e_2800;
    logic[7:0] _e_2801;
    (* src = "src/generated_driver.spade:846,2" *)
    logic[15:0] _e_2799;
    logic[7:0] _e_2803;
    logic[7:0] _e_2804;
    (* src = "src/generated_driver.spade:847,2" *)
    logic[15:0] _e_2802;
    logic[7:0] _e_2806;
    logic[7:0] _e_2807;
    (* src = "src/generated_driver.spade:848,2" *)
    logic[15:0] _e_2805;
    logic[7:0] _e_2809;
    logic[7:0] _e_2810;
    (* src = "src/generated_driver.spade:849,2" *)
    logic[15:0] _e_2808;
    logic[7:0] _e_2812;
    logic[7:0] _e_2813;
    (* src = "src/generated_driver.spade:850,2" *)
    logic[15:0] _e_2811;
    logic[7:0] _e_2815;
    logic[7:0] _e_2816;
    (* src = "src/generated_driver.spade:851,2" *)
    logic[15:0] _e_2814;
    logic[7:0] _e_2818;
    logic[7:0] _e_2819;
    (* src = "src/generated_driver.spade:852,2" *)
    logic[15:0] _e_2817;
    logic[7:0] _e_2821;
    logic[7:0] _e_2822;
    (* src = "src/generated_driver.spade:853,2" *)
    logic[15:0] _e_2820;
    logic[7:0] _e_2824;
    logic[7:0] _e_2825;
    (* src = "src/generated_driver.spade:854,2" *)
    logic[15:0] _e_2823;
    logic[7:0] _e_2827;
    logic[7:0] _e_2828;
    (* src = "src/generated_driver.spade:855,2" *)
    logic[15:0] _e_2826;
    logic[7:0] _e_2830;
    logic[7:0] _e_2831;
    (* src = "src/generated_driver.spade:856,2" *)
    logic[15:0] _e_2829;
    logic[7:0] _e_2833;
    logic[7:0] _e_2834;
    (* src = "src/generated_driver.spade:857,2" *)
    logic[15:0] _e_2832;
    logic[7:0] _e_2836;
    logic[7:0] _e_2837;
    (* src = "src/generated_driver.spade:858,2" *)
    logic[15:0] _e_2835;
    logic[7:0] _e_2839;
    logic[7:0] _e_2840;
    (* src = "src/generated_driver.spade:859,2" *)
    logic[15:0] _e_2838;
    logic[7:0] _e_2842;
    logic[7:0] _e_2843;
    (* src = "src/generated_driver.spade:860,2" *)
    logic[15:0] _e_2841;
    logic[7:0] _e_2845;
    logic[7:0] _e_2846;
    (* src = "src/generated_driver.spade:861,2" *)
    logic[15:0] _e_2844;
    logic[7:0] _e_2848;
    logic[7:0] _e_2849;
    (* src = "src/generated_driver.spade:862,2" *)
    logic[15:0] _e_2847;
    logic[7:0] _e_2851;
    logic[7:0] _e_2852;
    (* src = "src/generated_driver.spade:863,2" *)
    logic[15:0] _e_2850;
    logic[7:0] _e_2854;
    logic[7:0] _e_2855;
    (* src = "src/generated_driver.spade:864,2" *)
    logic[15:0] _e_2853;
    logic[7:0] _e_2857;
    logic[7:0] _e_2858;
    (* src = "src/generated_driver.spade:865,2" *)
    logic[15:0] _e_2856;
    logic[7:0] _e_2860;
    logic[7:0] _e_2861;
    (* src = "src/generated_driver.spade:866,2" *)
    logic[15:0] _e_2859;
    logic[7:0] _e_2863;
    logic[7:0] _e_2864;
    (* src = "src/generated_driver.spade:867,2" *)
    logic[15:0] _e_2862;
    logic[7:0] _e_2866;
    logic[7:0] _e_2867;
    (* src = "src/generated_driver.spade:868,2" *)
    logic[15:0] _e_2865;
    logic[7:0] _e_2869;
    logic[7:0] _e_2870;
    (* src = "src/generated_driver.spade:869,2" *)
    logic[15:0] _e_2868;
    logic[7:0] _e_2872;
    logic[7:0] _e_2873;
    (* src = "src/generated_driver.spade:870,2" *)
    logic[15:0] _e_2871;
    logic[7:0] _e_2875;
    logic[7:0] _e_2876;
    (* src = "src/generated_driver.spade:871,2" *)
    logic[15:0] _e_2874;
    logic[7:0] _e_2878;
    logic[7:0] _e_2879;
    (* src = "src/generated_driver.spade:872,2" *)
    logic[15:0] _e_2877;
    logic[7:0] _e_2881;
    logic[7:0] _e_2882;
    (* src = "src/generated_driver.spade:873,2" *)
    logic[15:0] _e_2880;
    logic[7:0] _e_2884;
    logic[7:0] _e_2885;
    (* src = "src/generated_driver.spade:874,2" *)
    logic[15:0] _e_2883;
    logic[7:0] _e_2887;
    logic[7:0] _e_2888;
    (* src = "src/generated_driver.spade:875,2" *)
    logic[15:0] _e_2886;
    logic[7:0] _e_2890;
    logic[7:0] _e_2891;
    (* src = "src/generated_driver.spade:876,2" *)
    logic[15:0] _e_2889;
    logic[7:0] _e_2893;
    logic[7:0] _e_2894;
    (* src = "src/generated_driver.spade:877,2" *)
    logic[15:0] _e_2892;
    logic[7:0] _e_2896;
    logic[7:0] _e_2897;
    (* src = "src/generated_driver.spade:878,2" *)
    logic[15:0] _e_2895;
    logic[7:0] _e_2899;
    logic[7:0] _e_2900;
    (* src = "src/generated_driver.spade:879,2" *)
    logic[15:0] _e_2898;
    logic[7:0] _e_2902;
    logic[7:0] _e_2903;
    (* src = "src/generated_driver.spade:880,2" *)
    logic[15:0] _e_2901;
    logic[7:0] _e_2905;
    logic[7:0] _e_2906;
    (* src = "src/generated_driver.spade:881,2" *)
    logic[15:0] _e_2904;
    logic[7:0] _e_2908;
    logic[7:0] _e_2909;
    (* src = "src/generated_driver.spade:882,2" *)
    logic[15:0] _e_2907;
    logic[7:0] _e_2911;
    logic[7:0] _e_2912;
    (* src = "src/generated_driver.spade:883,2" *)
    logic[15:0] _e_2910;
    logic[7:0] _e_2914;
    logic[7:0] _e_2915;
    (* src = "src/generated_driver.spade:884,2" *)
    logic[15:0] _e_2913;
    logic[7:0] _e_2917;
    logic[7:0] _e_2918;
    (* src = "src/generated_driver.spade:885,2" *)
    logic[15:0] _e_2916;
    logic[7:0] _e_2920;
    logic[7:0] _e_2921;
    (* src = "src/generated_driver.spade:886,2" *)
    logic[15:0] _e_2919;
    logic[7:0] _e_2923;
    logic[7:0] _e_2924;
    (* src = "src/generated_driver.spade:887,2" *)
    logic[15:0] _e_2922;
    logic[7:0] _e_2926;
    logic[7:0] _e_2927;
    (* src = "src/generated_driver.spade:888,2" *)
    logic[15:0] _e_2925;
    logic[7:0] _e_2929;
    logic[7:0] _e_2930;
    (* src = "src/generated_driver.spade:889,2" *)
    logic[15:0] _e_2928;
    logic[7:0] _e_2932;
    logic[7:0] _e_2933;
    (* src = "src/generated_driver.spade:890,2" *)
    logic[15:0] _e_2931;
    logic[7:0] _e_2935;
    logic[7:0] _e_2936;
    (* src = "src/generated_driver.spade:891,2" *)
    logic[15:0] _e_2934;
    logic[7:0] _e_2938;
    logic[7:0] _e_2939;
    (* src = "src/generated_driver.spade:892,2" *)
    logic[15:0] _e_2937;
    logic[7:0] _e_2941;
    logic[7:0] _e_2942;
    (* src = "src/generated_driver.spade:893,2" *)
    logic[15:0] _e_2940;
    logic[7:0] _e_2944;
    logic[7:0] _e_2945;
    (* src = "src/generated_driver.spade:894,2" *)
    logic[15:0] _e_2943;
    logic[7:0] _e_2947;
    logic[7:0] _e_2948;
    (* src = "src/generated_driver.spade:895,2" *)
    logic[15:0] _e_2946;
    logic[7:0] _e_2950;
    logic[7:0] _e_2951;
    (* src = "src/generated_driver.spade:896,2" *)
    logic[15:0] _e_2949;
    logic[7:0] _e_2953;
    logic[7:0] _e_2954;
    (* src = "src/generated_driver.spade:897,2" *)
    logic[15:0] _e_2952;
    logic[7:0] _e_2956;
    logic[7:0] _e_2957;
    (* src = "src/generated_driver.spade:898,2" *)
    logic[15:0] _e_2955;
    logic[7:0] _e_2959;
    logic[7:0] _e_2960;
    (* src = "src/generated_driver.spade:899,2" *)
    logic[15:0] _e_2958;
    logic[7:0] _e_2962;
    logic[7:0] _e_2963;
    (* src = "src/generated_driver.spade:900,2" *)
    logic[15:0] _e_2961;
    logic[7:0] _e_2965;
    logic[7:0] _e_2966;
    (* src = "src/generated_driver.spade:901,2" *)
    logic[15:0] _e_2964;
    logic[7:0] _e_2968;
    logic[7:0] _e_2969;
    (* src = "src/generated_driver.spade:902,2" *)
    logic[15:0] _e_2967;
    logic[7:0] _e_2971;
    logic[7:0] _e_2972;
    (* src = "src/generated_driver.spade:903,2" *)
    logic[15:0] _e_2970;
    logic[7:0] _e_2974;
    logic[7:0] _e_2975;
    (* src = "src/generated_driver.spade:904,2" *)
    logic[15:0] _e_2973;
    logic[7:0] _e_2977;
    logic[7:0] _e_2978;
    (* src = "src/generated_driver.spade:905,2" *)
    logic[15:0] _e_2976;
    logic[7:0] _e_2980;
    logic[7:0] _e_2981;
    (* src = "src/generated_driver.spade:906,2" *)
    logic[15:0] _e_2979;
    logic[7:0] _e_2983;
    logic[7:0] _e_2984;
    (* src = "src/generated_driver.spade:907,2" *)
    logic[15:0] _e_2982;
    logic[7:0] _e_2986;
    logic[7:0] _e_2987;
    (* src = "src/generated_driver.spade:908,2" *)
    logic[15:0] _e_2985;
    logic[7:0] _e_2989;
    logic[7:0] _e_2990;
    (* src = "src/generated_driver.spade:909,2" *)
    logic[15:0] _e_2988;
    logic[7:0] _e_2992;
    logic[7:0] _e_2993;
    (* src = "src/generated_driver.spade:910,2" *)
    logic[15:0] _e_2991;
    logic[7:0] _e_2995;
    logic[7:0] _e_2996;
    (* src = "src/generated_driver.spade:911,2" *)
    logic[15:0] _e_2994;
    logic[7:0] _e_2998;
    logic[7:0] _e_2999;
    (* src = "src/generated_driver.spade:912,2" *)
    logic[15:0] _e_2997;
    logic[7:0] _e_3001;
    logic[7:0] _e_3002;
    (* src = "src/generated_driver.spade:913,2" *)
    logic[15:0] _e_3000;
    logic[7:0] _e_3004;
    logic[7:0] _e_3005;
    (* src = "src/generated_driver.spade:914,2" *)
    logic[15:0] _e_3003;
    logic[7:0] _e_3007;
    logic[7:0] _e_3008;
    (* src = "src/generated_driver.spade:915,2" *)
    logic[15:0] _e_3006;
    logic[7:0] _e_3010;
    logic[7:0] _e_3011;
    (* src = "src/generated_driver.spade:916,2" *)
    logic[15:0] _e_3009;
    logic[7:0] _e_3013;
    logic[7:0] _e_3014;
    (* src = "src/generated_driver.spade:917,2" *)
    logic[15:0] _e_3012;
    logic[7:0] _e_3016;
    logic[7:0] _e_3017;
    (* src = "src/generated_driver.spade:918,2" *)
    logic[15:0] _e_3015;
    logic[7:0] _e_3019;
    logic[7:0] _e_3020;
    (* src = "src/generated_driver.spade:919,2" *)
    logic[15:0] _e_3018;
    logic[7:0] _e_3022;
    logic[7:0] _e_3023;
    (* src = "src/generated_driver.spade:920,2" *)
    logic[15:0] _e_3021;
    logic[7:0] _e_3025;
    logic[7:0] _e_3026;
    (* src = "src/generated_driver.spade:921,2" *)
    logic[15:0] _e_3024;
    logic[7:0] _e_3028;
    logic[7:0] _e_3029;
    (* src = "src/generated_driver.spade:922,2" *)
    logic[15:0] _e_3027;
    logic[7:0] _e_3031;
    logic[7:0] _e_3032;
    (* src = "src/generated_driver.spade:923,2" *)
    logic[15:0] _e_3030;
    logic[7:0] _e_3034;
    logic[7:0] _e_3035;
    (* src = "src/generated_driver.spade:924,2" *)
    logic[15:0] _e_3033;
    logic[7:0] _e_3037;
    logic[7:0] _e_3038;
    (* src = "src/generated_driver.spade:925,2" *)
    logic[15:0] _e_3036;
    logic[7:0] _e_3040;
    logic[7:0] _e_3041;
    (* src = "src/generated_driver.spade:926,2" *)
    logic[15:0] _e_3039;
    logic[7:0] _e_3043;
    logic[7:0] _e_3044;
    (* src = "src/generated_driver.spade:927,2" *)
    logic[15:0] _e_3042;
    logic[7:0] _e_3046;
    logic[7:0] _e_3047;
    (* src = "src/generated_driver.spade:928,2" *)
    logic[15:0] _e_3045;
    logic[7:0] _e_3049;
    logic[7:0] _e_3050;
    (* src = "src/generated_driver.spade:929,2" *)
    logic[15:0] _e_3048;
    logic[7:0] _e_3052;
    logic[7:0] _e_3053;
    (* src = "src/generated_driver.spade:930,2" *)
    logic[15:0] _e_3051;
    logic[7:0] _e_3055;
    logic[7:0] _e_3056;
    (* src = "src/generated_driver.spade:931,2" *)
    logic[15:0] _e_3054;
    logic[7:0] _e_3058;
    logic[7:0] _e_3059;
    (* src = "src/generated_driver.spade:932,2" *)
    logic[15:0] _e_3057;
    logic[7:0] _e_3061;
    logic[7:0] _e_3062;
    (* src = "src/generated_driver.spade:933,2" *)
    logic[15:0] _e_3060;
    logic[7:0] _e_3064;
    logic[7:0] _e_3065;
    (* src = "src/generated_driver.spade:934,2" *)
    logic[15:0] _e_3063;
    logic[7:0] _e_3067;
    logic[7:0] _e_3068;
    (* src = "src/generated_driver.spade:935,2" *)
    logic[15:0] _e_3066;
    logic[7:0] _e_3070;
    logic[7:0] _e_3071;
    (* src = "src/generated_driver.spade:936,2" *)
    logic[15:0] _e_3069;
    logic[7:0] _e_3073;
    logic[7:0] _e_3074;
    (* src = "src/generated_driver.spade:937,2" *)
    logic[15:0] _e_3072;
    logic[7:0] _e_3076;
    logic[7:0] _e_3077;
    (* src = "src/generated_driver.spade:938,2" *)
    logic[15:0] _e_3075;
    logic[7:0] _e_3079;
    logic[7:0] _e_3080;
    (* src = "src/generated_driver.spade:939,2" *)
    logic[15:0] _e_3078;
    logic[7:0] _e_3082;
    logic[7:0] _e_3083;
    (* src = "src/generated_driver.spade:940,2" *)
    logic[15:0] _e_3081;
    logic[7:0] _e_3085;
    logic[7:0] _e_3086;
    (* src = "src/generated_driver.spade:941,2" *)
    logic[15:0] _e_3084;
    logic[7:0] _e_3088;
    logic[7:0] _e_3089;
    (* src = "src/generated_driver.spade:942,2" *)
    logic[15:0] _e_3087;
    logic[7:0] _e_3091;
    logic[7:0] _e_3092;
    (* src = "src/generated_driver.spade:943,2" *)
    logic[15:0] _e_3090;
    logic[7:0] _e_3094;
    logic[7:0] _e_3095;
    (* src = "src/generated_driver.spade:944,2" *)
    logic[15:0] _e_3093;
    logic[7:0] _e_3097;
    logic[7:0] _e_3098;
    (* src = "src/generated_driver.spade:945,2" *)
    logic[15:0] _e_3096;
    logic[7:0] _e_3100;
    logic[7:0] _e_3101;
    (* src = "src/generated_driver.spade:946,2" *)
    logic[15:0] _e_3099;
    logic[7:0] _e_3103;
    logic[7:0] _e_3104;
    (* src = "src/generated_driver.spade:947,2" *)
    logic[15:0] _e_3102;
    logic[7:0] _e_3106;
    logic[7:0] _e_3107;
    (* src = "src/generated_driver.spade:948,2" *)
    logic[15:0] _e_3105;
    logic[7:0] _e_3109;
    logic[7:0] _e_3110;
    (* src = "src/generated_driver.spade:949,2" *)
    logic[15:0] _e_3108;
    logic[7:0] _e_3112;
    logic[7:0] _e_3113;
    (* src = "src/generated_driver.spade:950,2" *)
    logic[15:0] _e_3111;
    logic[7:0] _e_3115;
    logic[7:0] _e_3116;
    (* src = "src/generated_driver.spade:951,2" *)
    logic[15:0] _e_3114;
    logic[7:0] _e_3118;
    logic[7:0] _e_3119;
    (* src = "src/generated_driver.spade:952,2" *)
    logic[15:0] _e_3117;
    logic[7:0] _e_3121;
    logic[7:0] _e_3122;
    (* src = "src/generated_driver.spade:953,2" *)
    logic[15:0] _e_3120;
    logic[7:0] _e_3124;
    logic[7:0] _e_3125;
    (* src = "src/generated_driver.spade:954,2" *)
    logic[15:0] _e_3123;
    logic[7:0] _e_3127;
    logic[7:0] _e_3128;
    (* src = "src/generated_driver.spade:955,2" *)
    logic[15:0] _e_3126;
    logic[7:0] _e_3130;
    logic[7:0] _e_3131;
    (* src = "src/generated_driver.spade:956,2" *)
    logic[15:0] _e_3129;
    logic[7:0] _e_3133;
    logic[7:0] _e_3134;
    (* src = "src/generated_driver.spade:957,2" *)
    logic[15:0] _e_3132;
    logic[7:0] _e_3136;
    logic[7:0] _e_3137;
    (* src = "src/generated_driver.spade:958,2" *)
    logic[15:0] _e_3135;
    logic[7:0] _e_3139;
    logic[7:0] _e_3140;
    (* src = "src/generated_driver.spade:959,2" *)
    logic[15:0] _e_3138;
    logic[7:0] _e_3142;
    logic[7:0] _e_3143;
    (* src = "src/generated_driver.spade:960,2" *)
    logic[15:0] _e_3141;
    logic[7:0] _e_3145;
    logic[7:0] _e_3146;
    (* src = "src/generated_driver.spade:961,2" *)
    logic[15:0] _e_3144;
    logic[7:0] _e_3148;
    logic[7:0] _e_3149;
    (* src = "src/generated_driver.spade:962,2" *)
    logic[15:0] _e_3147;
    logic[7:0] _e_3151;
    logic[7:0] _e_3152;
    (* src = "src/generated_driver.spade:963,2" *)
    logic[15:0] _e_3150;
    logic[7:0] _e_3154;
    logic[7:0] _e_3155;
    (* src = "src/generated_driver.spade:964,2" *)
    logic[15:0] _e_3153;
    logic[7:0] _e_3157;
    logic[7:0] _e_3158;
    (* src = "src/generated_driver.spade:965,2" *)
    logic[15:0] _e_3156;
    logic[7:0] _e_3160;
    logic[7:0] _e_3161;
    (* src = "src/generated_driver.spade:966,2" *)
    logic[15:0] _e_3159;
    logic[7:0] _e_3163;
    logic[7:0] _e_3164;
    (* src = "src/generated_driver.spade:967,2" *)
    logic[15:0] _e_3162;
    logic[7:0] _e_3166;
    logic[7:0] _e_3167;
    (* src = "src/generated_driver.spade:968,2" *)
    logic[15:0] _e_3165;
    logic[7:0] _e_3169;
    logic[7:0] _e_3170;
    (* src = "src/generated_driver.spade:969,2" *)
    logic[15:0] _e_3168;
    logic[7:0] _e_3172;
    logic[7:0] _e_3173;
    (* src = "src/generated_driver.spade:970,2" *)
    logic[15:0] _e_3171;
    logic[7:0] _e_3175;
    logic[7:0] _e_3176;
    (* src = "src/generated_driver.spade:971,2" *)
    logic[15:0] _e_3174;
    logic[7:0] _e_3178;
    logic[7:0] _e_3179;
    (* src = "src/generated_driver.spade:972,2" *)
    logic[15:0] _e_3177;
    logic[7:0] _e_3181;
    logic[7:0] _e_3182;
    (* src = "src/generated_driver.spade:973,2" *)
    logic[15:0] _e_3180;
    logic[7:0] _e_3184;
    logic[7:0] _e_3185;
    (* src = "src/generated_driver.spade:974,2" *)
    logic[15:0] _e_3183;
    logic[7:0] _e_3187;
    logic[7:0] _e_3188;
    (* src = "src/generated_driver.spade:975,2" *)
    logic[15:0] _e_3186;
    logic[7:0] _e_3190;
    logic[7:0] _e_3191;
    (* src = "src/generated_driver.spade:976,2" *)
    logic[15:0] _e_3189;
    logic[7:0] _e_3193;
    logic[7:0] _e_3194;
    (* src = "src/generated_driver.spade:977,2" *)
    logic[15:0] _e_3192;
    logic[7:0] _e_3196;
    logic[7:0] _e_3197;
    (* src = "src/generated_driver.spade:978,2" *)
    logic[15:0] _e_3195;
    logic[7:0] _e_3199;
    logic[7:0] _e_3200;
    (* src = "src/generated_driver.spade:979,2" *)
    logic[15:0] _e_3198;
    logic[7:0] _e_3202;
    logic[7:0] _e_3203;
    (* src = "src/generated_driver.spade:980,2" *)
    logic[15:0] _e_3201;
    logic[7:0] _e_3205;
    logic[7:0] _e_3206;
    (* src = "src/generated_driver.spade:981,2" *)
    logic[15:0] _e_3204;
    logic[7:0] _e_3208;
    logic[7:0] _e_3209;
    (* src = "src/generated_driver.spade:982,2" *)
    logic[15:0] _e_3207;
    logic[7:0] _e_3211;
    logic[7:0] _e_3212;
    (* src = "src/generated_driver.spade:983,2" *)
    logic[15:0] _e_3210;
    logic[7:0] _e_3214;
    logic[7:0] _e_3215;
    (* src = "src/generated_driver.spade:984,2" *)
    logic[15:0] _e_3213;
    logic[7:0] _e_3217;
    logic[7:0] _e_3218;
    (* src = "src/generated_driver.spade:985,2" *)
    logic[15:0] _e_3216;
    logic[7:0] _e_3220;
    logic[7:0] _e_3221;
    (* src = "src/generated_driver.spade:986,2" *)
    logic[15:0] _e_3219;
    logic[7:0] _e_3223;
    logic[7:0] _e_3224;
    (* src = "src/generated_driver.spade:987,2" *)
    logic[15:0] _e_3222;
    logic[7:0] _e_3226;
    logic[7:0] _e_3227;
    (* src = "src/generated_driver.spade:988,2" *)
    logic[15:0] _e_3225;
    logic[7:0] _e_3229;
    logic[7:0] _e_3230;
    (* src = "src/generated_driver.spade:989,2" *)
    logic[15:0] _e_3228;
    logic[7:0] _e_3232;
    logic[7:0] _e_3233;
    (* src = "src/generated_driver.spade:990,2" *)
    logic[15:0] _e_3231;
    logic[7:0] _e_3235;
    logic[7:0] _e_3236;
    (* src = "src/generated_driver.spade:991,2" *)
    logic[15:0] _e_3234;
    logic[7:0] _e_3238;
    logic[7:0] _e_3239;
    (* src = "src/generated_driver.spade:992,2" *)
    logic[15:0] _e_3237;
    logic[7:0] _e_3241;
    logic[7:0] _e_3242;
    (* src = "src/generated_driver.spade:993,2" *)
    logic[15:0] _e_3240;
    logic[7:0] _e_3244;
    logic[7:0] _e_3245;
    (* src = "src/generated_driver.spade:994,2" *)
    logic[15:0] _e_3243;
    logic[7:0] _e_3247;
    logic[7:0] _e_3248;
    (* src = "src/generated_driver.spade:995,2" *)
    logic[15:0] _e_3246;
    logic[7:0] _e_3250;
    logic[7:0] _e_3251;
    (* src = "src/generated_driver.spade:996,2" *)
    logic[15:0] _e_3249;
    logic[7:0] _e_3253;
    logic[7:0] _e_3254;
    (* src = "src/generated_driver.spade:997,2" *)
    logic[15:0] _e_3252;
    logic[7:0] _e_3256;
    logic[7:0] _e_3257;
    (* src = "src/generated_driver.spade:998,2" *)
    logic[15:0] _e_3255;
    logic[7:0] _e_3259;
    logic[7:0] _e_3260;
    (* src = "src/generated_driver.spade:999,2" *)
    logic[15:0] _e_3258;
    logic[7:0] _e_3262;
    logic[7:0] _e_3263;
    (* src = "src/generated_driver.spade:1000,2" *)
    logic[15:0] _e_3261;
    logic[7:0] _e_3265;
    logic[7:0] _e_3266;
    (* src = "src/generated_driver.spade:1001,2" *)
    logic[15:0] _e_3264;
    logic[7:0] _e_3268;
    logic[7:0] _e_3269;
    (* src = "src/generated_driver.spade:1002,2" *)
    logic[15:0] _e_3267;
    logic[7:0] _e_3271;
    logic[7:0] _e_3272;
    (* src = "src/generated_driver.spade:1003,2" *)
    logic[15:0] _e_3270;
    logic[7:0] _e_3274;
    logic[7:0] _e_3275;
    (* src = "src/generated_driver.spade:1004,2" *)
    logic[15:0] _e_3273;
    logic[7:0] _e_3277;
    logic[7:0] _e_3278;
    (* src = "src/generated_driver.spade:1005,2" *)
    logic[15:0] _e_3276;
    logic[7:0] _e_3280;
    logic[7:0] _e_3281;
    (* src = "src/generated_driver.spade:1006,2" *)
    logic[15:0] _e_3279;
    logic[7:0] _e_3283;
    logic[7:0] _e_3284;
    (* src = "src/generated_driver.spade:1007,2" *)
    logic[15:0] _e_3282;
    logic[7:0] _e_3286;
    logic[7:0] _e_3287;
    (* src = "src/generated_driver.spade:1008,2" *)
    logic[15:0] _e_3285;
    logic[7:0] _e_3289;
    logic[7:0] _e_3290;
    (* src = "src/generated_driver.spade:1009,2" *)
    logic[15:0] _e_3288;
    logic[7:0] _e_3292;
    logic[7:0] _e_3293;
    (* src = "src/generated_driver.spade:1010,2" *)
    logic[15:0] _e_3291;
    logic[7:0] _e_3295;
    logic[7:0] _e_3296;
    (* src = "src/generated_driver.spade:1011,2" *)
    logic[15:0] _e_3294;
    logic[7:0] _e_3298;
    logic[7:0] _e_3299;
    (* src = "src/generated_driver.spade:1012,2" *)
    logic[15:0] _e_3297;
    logic[7:0] _e_3301;
    logic[7:0] _e_3302;
    (* src = "src/generated_driver.spade:1013,2" *)
    logic[15:0] _e_3300;
    logic[7:0] _e_3304;
    logic[7:0] _e_3305;
    (* src = "src/generated_driver.spade:1014,2" *)
    logic[15:0] _e_3303;
    logic[7:0] _e_3307;
    logic[7:0] _e_3308;
    (* src = "src/generated_driver.spade:1015,2" *)
    logic[15:0] _e_3306;
    logic[7:0] _e_3310;
    logic[7:0] _e_3311;
    (* src = "src/generated_driver.spade:1016,2" *)
    logic[15:0] _e_3309;
    logic[7:0] _e_3313;
    logic[7:0] _e_3314;
    (* src = "src/generated_driver.spade:1017,2" *)
    logic[15:0] _e_3312;
    logic[7:0] _e_3316;
    logic[7:0] _e_3317;
    (* src = "src/generated_driver.spade:1018,2" *)
    logic[15:0] _e_3315;
    logic[7:0] _e_3319;
    logic[7:0] _e_3320;
    (* src = "src/generated_driver.spade:1019,2" *)
    logic[15:0] _e_3318;
    logic[7:0] _e_3322;
    logic[7:0] _e_3323;
    (* src = "src/generated_driver.spade:1020,2" *)
    logic[15:0] _e_3321;
    logic[7:0] _e_3325;
    logic[7:0] _e_3326;
    (* src = "src/generated_driver.spade:1021,2" *)
    logic[15:0] _e_3324;
    logic[7:0] _e_3328;
    logic[7:0] _e_3329;
    (* src = "src/generated_driver.spade:1022,2" *)
    logic[15:0] _e_3327;
    logic[7:0] _e_3331;
    logic[7:0] _e_3332;
    (* src = "src/generated_driver.spade:1023,2" *)
    logic[15:0] _e_3330;
    logic[7:0] _e_3334;
    logic[7:0] _e_3335;
    (* src = "src/generated_driver.spade:1024,2" *)
    logic[15:0] _e_3333;
    logic[7:0] _e_3337;
    logic[7:0] _e_3338;
    (* src = "src/generated_driver.spade:1025,2" *)
    logic[15:0] _e_3336;
    logic[7:0] _e_3340;
    logic[7:0] _e_3341;
    (* src = "src/generated_driver.spade:1026,2" *)
    logic[15:0] _e_3339;
    logic[7:0] _e_3343;
    logic[7:0] _e_3344;
    (* src = "src/generated_driver.spade:1027,2" *)
    logic[15:0] _e_3342;
    logic[7:0] _e_3346;
    logic[7:0] _e_3347;
    (* src = "src/generated_driver.spade:1028,2" *)
    logic[15:0] _e_3345;
    logic[7:0] _e_3349;
    logic[7:0] _e_3350;
    (* src = "src/generated_driver.spade:1029,2" *)
    logic[15:0] _e_3348;
    logic[7:0] _e_3352;
    logic[7:0] _e_3353;
    (* src = "src/generated_driver.spade:1030,2" *)
    logic[15:0] _e_3351;
    logic[7:0] _e_3355;
    logic[7:0] _e_3356;
    (* src = "src/generated_driver.spade:1031,2" *)
    logic[15:0] _e_3354;
    logic[7:0] _e_3358;
    logic[7:0] _e_3359;
    (* src = "src/generated_driver.spade:1032,2" *)
    logic[15:0] _e_3357;
    logic[7:0] _e_3361;
    logic[7:0] _e_3362;
    (* src = "src/generated_driver.spade:1033,2" *)
    logic[15:0] _e_3360;
    logic[7:0] _e_3364;
    logic[7:0] _e_3365;
    (* src = "src/generated_driver.spade:1034,2" *)
    logic[15:0] _e_3363;
    logic[7:0] _e_3367;
    logic[7:0] _e_3368;
    (* src = "src/generated_driver.spade:1035,2" *)
    logic[15:0] _e_3366;
    logic[7:0] _e_3370;
    logic[7:0] _e_3371;
    (* src = "src/generated_driver.spade:1036,2" *)
    logic[15:0] _e_3369;
    logic[7:0] _e_3373;
    logic[7:0] _e_3374;
    (* src = "src/generated_driver.spade:1037,2" *)
    logic[15:0] _e_3372;
    logic[7:0] _e_3376;
    logic[7:0] _e_3377;
    (* src = "src/generated_driver.spade:1038,2" *)
    logic[15:0] _e_3375;
    logic[7:0] _e_3379;
    logic[7:0] _e_3380;
    (* src = "src/generated_driver.spade:1039,2" *)
    logic[15:0] _e_3378;
    logic[7:0] _e_3382;
    logic[7:0] _e_3383;
    (* src = "src/generated_driver.spade:1040,2" *)
    logic[15:0] _e_3381;
    logic[7:0] _e_3385;
    logic[7:0] _e_3386;
    (* src = "src/generated_driver.spade:1041,2" *)
    logic[15:0] _e_3384;
    logic[7:0] _e_3388;
    logic[7:0] _e_3389;
    (* src = "src/generated_driver.spade:1042,2" *)
    logic[15:0] _e_3387;
    logic[7:0] _e_3391;
    logic[7:0] _e_3392;
    (* src = "src/generated_driver.spade:1043,2" *)
    logic[15:0] _e_3390;
    logic[7:0] _e_3394;
    logic[7:0] _e_3395;
    (* src = "src/generated_driver.spade:1044,2" *)
    logic[15:0] _e_3393;
    logic[7:0] _e_3397;
    logic[7:0] _e_3398;
    (* src = "src/generated_driver.spade:1045,2" *)
    logic[15:0] _e_3396;
    logic[7:0] _e_3400;
    logic[7:0] _e_3401;
    (* src = "src/generated_driver.spade:1046,2" *)
    logic[15:0] _e_3399;
    logic[7:0] _e_3403;
    logic[7:0] _e_3404;
    (* src = "src/generated_driver.spade:1047,2" *)
    logic[15:0] _e_3402;
    logic[7:0] _e_3406;
    logic[7:0] _e_3407;
    (* src = "src/generated_driver.spade:1048,2" *)
    logic[15:0] _e_3405;
    logic[7:0] _e_3409;
    logic[7:0] _e_3410;
    (* src = "src/generated_driver.spade:1049,2" *)
    logic[15:0] _e_3408;
    logic[7:0] _e_3412;
    logic[7:0] _e_3413;
    (* src = "src/generated_driver.spade:1050,2" *)
    logic[15:0] _e_3411;
    logic[7:0] _e_3415;
    logic[7:0] _e_3416;
    (* src = "src/generated_driver.spade:1051,2" *)
    logic[15:0] _e_3414;
    logic[7:0] _e_3418;
    logic[7:0] _e_3419;
    (* src = "src/generated_driver.spade:1052,2" *)
    logic[15:0] _e_3417;
    logic[7:0] _e_3421;
    logic[7:0] _e_3422;
    (* src = "src/generated_driver.spade:1053,2" *)
    logic[15:0] _e_3420;
    logic[7:0] _e_3424;
    logic[7:0] _e_3425;
    (* src = "src/generated_driver.spade:1054,2" *)
    logic[15:0] _e_3423;
    logic[7:0] _e_3427;
    logic[7:0] _e_3428;
    (* src = "src/generated_driver.spade:1055,2" *)
    logic[15:0] _e_3426;
    logic[7:0] _e_3430;
    logic[7:0] _e_3431;
    (* src = "src/generated_driver.spade:1056,2" *)
    logic[15:0] _e_3429;
    logic[7:0] _e_3433;
    logic[7:0] _e_3434;
    (* src = "src/generated_driver.spade:1057,2" *)
    logic[15:0] _e_3432;
    logic[7:0] _e_3436;
    logic[7:0] _e_3437;
    (* src = "src/generated_driver.spade:1058,2" *)
    logic[15:0] _e_3435;
    logic[7:0] _e_3439;
    logic[7:0] _e_3440;
    (* src = "src/generated_driver.spade:1059,2" *)
    logic[15:0] _e_3438;
    logic[7:0] _e_3442;
    logic[7:0] _e_3443;
    (* src = "src/generated_driver.spade:1060,2" *)
    logic[15:0] _e_3441;
    logic[7:0] _e_3445;
    logic[7:0] _e_3446;
    (* src = "src/generated_driver.spade:1061,2" *)
    logic[15:0] _e_3444;
    logic[7:0] _e_3448;
    logic[7:0] _e_3449;
    (* src = "src/generated_driver.spade:1062,2" *)
    logic[15:0] _e_3447;
    logic[7:0] _e_3451;
    logic[7:0] _e_3452;
    (* src = "src/generated_driver.spade:1063,2" *)
    logic[15:0] _e_3450;
    logic[7:0] _e_3454;
    logic[7:0] _e_3455;
    (* src = "src/generated_driver.spade:1064,2" *)
    logic[15:0] _e_3453;
    logic[7:0] _e_3457;
    logic[7:0] _e_3458;
    (* src = "src/generated_driver.spade:1065,2" *)
    logic[15:0] _e_3456;
    logic[7:0] _e_3460;
    logic[7:0] _e_3461;
    (* src = "src/generated_driver.spade:1066,2" *)
    logic[15:0] _e_3459;
    logic[7:0] _e_3463;
    logic[7:0] _e_3464;
    (* src = "src/generated_driver.spade:1067,2" *)
    logic[15:0] _e_3462;
    logic[7:0] _e_3466;
    logic[7:0] _e_3467;
    (* src = "src/generated_driver.spade:1068,2" *)
    logic[15:0] _e_3465;
    logic[7:0] _e_3469;
    logic[7:0] _e_3470;
    (* src = "src/generated_driver.spade:1069,2" *)
    logic[15:0] _e_3468;
    logic[7:0] _e_3472;
    logic[7:0] _e_3473;
    (* src = "src/generated_driver.spade:1070,2" *)
    logic[15:0] _e_3471;
    logic[7:0] _e_3475;
    logic[7:0] _e_3476;
    (* src = "src/generated_driver.spade:1071,2" *)
    logic[15:0] _e_3474;
    logic[7:0] _e_3478;
    logic[7:0] _e_3479;
    (* src = "src/generated_driver.spade:1072,2" *)
    logic[15:0] _e_3477;
    logic[7:0] _e_3481;
    logic[7:0] _e_3482;
    (* src = "src/generated_driver.spade:1073,2" *)
    logic[15:0] _e_3480;
    logic[7:0] _e_3484;
    logic[7:0] _e_3485;
    (* src = "src/generated_driver.spade:1074,2" *)
    logic[15:0] _e_3483;
    logic[7:0] _e_3487;
    logic[7:0] _e_3488;
    (* src = "src/generated_driver.spade:1075,2" *)
    logic[15:0] _e_3486;
    logic[7:0] _e_3490;
    logic[7:0] _e_3491;
    (* src = "src/generated_driver.spade:1076,2" *)
    logic[15:0] _e_3489;
    logic[7:0] _e_3493;
    logic[7:0] _e_3494;
    (* src = "src/generated_driver.spade:1077,2" *)
    logic[15:0] _e_3492;
    logic[7:0] _e_3496;
    logic[7:0] _e_3497;
    (* src = "src/generated_driver.spade:1078,2" *)
    logic[15:0] _e_3495;
    logic[7:0] _e_3499;
    logic[7:0] _e_3500;
    (* src = "src/generated_driver.spade:1079,2" *)
    logic[15:0] _e_3498;
    logic[7:0] _e_3502;
    logic[7:0] _e_3503;
    (* src = "src/generated_driver.spade:1080,2" *)
    logic[15:0] _e_3501;
    logic[7:0] _e_3505;
    logic[7:0] _e_3506;
    (* src = "src/generated_driver.spade:1081,2" *)
    logic[15:0] _e_3504;
    logic[7:0] _e_3508;
    logic[7:0] _e_3509;
    (* src = "src/generated_driver.spade:1082,2" *)
    logic[15:0] _e_3507;
    logic[7:0] _e_3511;
    logic[7:0] _e_3512;
    (* src = "src/generated_driver.spade:1083,2" *)
    logic[15:0] _e_3510;
    logic[7:0] _e_3514;
    logic[7:0] _e_3515;
    (* src = "src/generated_driver.spade:1084,2" *)
    logic[15:0] _e_3513;
    logic[7:0] _e_3517;
    logic[7:0] _e_3518;
    (* src = "src/generated_driver.spade:1085,2" *)
    logic[15:0] _e_3516;
    logic[7:0] _e_3520;
    logic[7:0] _e_3521;
    (* src = "src/generated_driver.spade:1086,2" *)
    logic[15:0] _e_3519;
    logic[7:0] _e_3523;
    logic[7:0] _e_3524;
    (* src = "src/generated_driver.spade:1087,2" *)
    logic[15:0] _e_3522;
    logic[7:0] _e_3526;
    logic[7:0] _e_3527;
    (* src = "src/generated_driver.spade:1088,2" *)
    logic[15:0] _e_3525;
    logic[7:0] _e_3529;
    logic[7:0] _e_3530;
    (* src = "src/generated_driver.spade:1089,2" *)
    logic[15:0] _e_3528;
    logic[7:0] _e_3532;
    logic[7:0] _e_3533;
    (* src = "src/generated_driver.spade:1090,2" *)
    logic[15:0] _e_3531;
    logic[7:0] _e_3535;
    logic[7:0] _e_3536;
    (* src = "src/generated_driver.spade:1091,2" *)
    logic[15:0] _e_3534;
    logic[7:0] _e_3538;
    logic[7:0] _e_3539;
    (* src = "src/generated_driver.spade:1092,2" *)
    logic[15:0] _e_3537;
    logic[7:0] _e_3541;
    logic[7:0] _e_3542;
    (* src = "src/generated_driver.spade:1093,2" *)
    logic[15:0] _e_3540;
    logic[7:0] _e_3544;
    logic[7:0] _e_3545;
    (* src = "src/generated_driver.spade:1094,2" *)
    logic[15:0] _e_3543;
    logic[7:0] _e_3547;
    logic[7:0] _e_3548;
    (* src = "src/generated_driver.spade:1095,2" *)
    logic[15:0] _e_3546;
    logic[7:0] _e_3550;
    logic[7:0] _e_3551;
    (* src = "src/generated_driver.spade:1096,2" *)
    logic[15:0] _e_3549;
    logic[7:0] _e_3553;
    logic[7:0] _e_3554;
    (* src = "src/generated_driver.spade:1097,2" *)
    logic[15:0] _e_3552;
    logic[7:0] _e_3556;
    logic[7:0] _e_3557;
    (* src = "src/generated_driver.spade:1098,2" *)
    logic[15:0] _e_3555;
    logic[7:0] _e_3559;
    logic[7:0] _e_3560;
    (* src = "src/generated_driver.spade:1099,2" *)
    logic[15:0] _e_3558;
    logic[7:0] _e_3562;
    logic[7:0] _e_3563;
    (* src = "src/generated_driver.spade:1100,2" *)
    logic[15:0] _e_3561;
    logic[7:0] _e_3565;
    logic[7:0] _e_3566;
    (* src = "src/generated_driver.spade:1101,2" *)
    logic[15:0] _e_3564;
    logic[7:0] _e_3568;
    logic[7:0] _e_3569;
    (* src = "src/generated_driver.spade:1102,2" *)
    logic[15:0] _e_3567;
    logic[7:0] _e_3571;
    logic[7:0] _e_3572;
    (* src = "src/generated_driver.spade:1103,2" *)
    logic[15:0] _e_3570;
    logic[7:0] _e_3574;
    logic[7:0] _e_3575;
    (* src = "src/generated_driver.spade:1104,2" *)
    logic[15:0] _e_3573;
    logic[7:0] _e_3577;
    logic[7:0] _e_3578;
    (* src = "src/generated_driver.spade:1105,2" *)
    logic[15:0] _e_3576;
    logic[7:0] _e_3580;
    logic[7:0] _e_3581;
    (* src = "src/generated_driver.spade:1106,2" *)
    logic[15:0] _e_3579;
    logic[7:0] _e_3583;
    logic[7:0] _e_3584;
    (* src = "src/generated_driver.spade:1107,2" *)
    logic[15:0] _e_3582;
    logic[7:0] _e_3586;
    logic[7:0] _e_3587;
    (* src = "src/generated_driver.spade:1108,2" *)
    logic[15:0] _e_3585;
    logic[7:0] _e_3589;
    logic[7:0] _e_3590;
    (* src = "src/generated_driver.spade:1109,2" *)
    logic[15:0] _e_3588;
    logic[7:0] _e_3592;
    logic[7:0] _e_3593;
    (* src = "src/generated_driver.spade:1110,2" *)
    logic[15:0] _e_3591;
    logic[7:0] _e_3595;
    logic[7:0] _e_3596;
    (* src = "src/generated_driver.spade:1111,2" *)
    logic[15:0] _e_3594;
    logic[7:0] _e_3598;
    logic[7:0] _e_3599;
    (* src = "src/generated_driver.spade:1112,2" *)
    logic[15:0] _e_3597;
    logic[7:0] _e_3601;
    logic[7:0] _e_3602;
    (* src = "src/generated_driver.spade:1113,2" *)
    logic[15:0] _e_3600;
    logic[7:0] _e_3604;
    logic[7:0] _e_3605;
    (* src = "src/generated_driver.spade:1114,2" *)
    logic[15:0] _e_3603;
    logic[7:0] _e_3607;
    logic[7:0] _e_3608;
    (* src = "src/generated_driver.spade:1115,2" *)
    logic[15:0] _e_3606;
    logic[7:0] _e_3610;
    logic[7:0] _e_3611;
    (* src = "src/generated_driver.spade:1116,2" *)
    logic[15:0] _e_3609;
    logic[7:0] _e_3613;
    logic[7:0] _e_3614;
    (* src = "src/generated_driver.spade:1117,2" *)
    logic[15:0] _e_3612;
    logic[7:0] _e_3616;
    logic[7:0] _e_3617;
    (* src = "src/generated_driver.spade:1118,2" *)
    logic[15:0] _e_3615;
    logic[7:0] _e_3619;
    logic[7:0] _e_3620;
    (* src = "src/generated_driver.spade:1119,2" *)
    logic[15:0] _e_3618;
    logic[7:0] _e_3622;
    logic[7:0] _e_3623;
    (* src = "src/generated_driver.spade:1120,2" *)
    logic[15:0] _e_3621;
    logic[7:0] _e_3625;
    logic[7:0] _e_3626;
    (* src = "src/generated_driver.spade:1121,2" *)
    logic[15:0] _e_3624;
    logic[7:0] _e_3628;
    logic[7:0] _e_3629;
    (* src = "src/generated_driver.spade:1122,2" *)
    logic[15:0] _e_3627;
    logic[7:0] _e_3631;
    logic[7:0] _e_3632;
    (* src = "src/generated_driver.spade:1123,2" *)
    logic[15:0] _e_3630;
    logic[7:0] _e_3634;
    logic[7:0] _e_3635;
    (* src = "src/generated_driver.spade:1124,2" *)
    logic[15:0] _e_3633;
    logic[7:0] _e_3637;
    logic[7:0] _e_3638;
    (* src = "src/generated_driver.spade:1125,2" *)
    logic[15:0] _e_3636;
    logic[7:0] _e_3640;
    logic[7:0] _e_3641;
    (* src = "src/generated_driver.spade:1126,2" *)
    logic[15:0] _e_3639;
    logic[7:0] _e_3643;
    logic[7:0] _e_3644;
    (* src = "src/generated_driver.spade:1127,2" *)
    logic[15:0] _e_3642;
    logic[7:0] _e_3646;
    logic[7:0] _e_3647;
    (* src = "src/generated_driver.spade:1128,2" *)
    logic[15:0] _e_3645;
    logic[7:0] _e_3649;
    logic[7:0] _e_3650;
    (* src = "src/generated_driver.spade:1129,2" *)
    logic[15:0] _e_3648;
    logic[7:0] _e_3652;
    logic[7:0] _e_3653;
    (* src = "src/generated_driver.spade:1130,2" *)
    logic[15:0] _e_3651;
    logic[7:0] _e_3655;
    logic[7:0] _e_3656;
    (* src = "src/generated_driver.spade:1131,2" *)
    logic[15:0] _e_3654;
    logic[7:0] _e_3658;
    logic[7:0] _e_3659;
    (* src = "src/generated_driver.spade:1132,2" *)
    logic[15:0] _e_3657;
    logic[7:0] _e_3661;
    logic[7:0] _e_3662;
    (* src = "src/generated_driver.spade:1133,2" *)
    logic[15:0] _e_3660;
    logic[7:0] _e_3664;
    logic[7:0] _e_3665;
    (* src = "src/generated_driver.spade:1134,2" *)
    logic[15:0] _e_3663;
    logic[7:0] _e_3667;
    logic[7:0] _e_3668;
    (* src = "src/generated_driver.spade:1135,2" *)
    logic[15:0] _e_3666;
    logic[7:0] _e_3670;
    logic[7:0] _e_3671;
    (* src = "src/generated_driver.spade:1136,2" *)
    logic[15:0] _e_3669;
    logic[7:0] _e_3673;
    logic[7:0] _e_3674;
    (* src = "src/generated_driver.spade:1137,2" *)
    logic[15:0] _e_3672;
    logic[7:0] _e_3676;
    logic[7:0] _e_3677;
    (* src = "src/generated_driver.spade:1138,2" *)
    logic[15:0] _e_3675;
    logic[7:0] _e_3679;
    logic[7:0] _e_3680;
    (* src = "src/generated_driver.spade:1139,2" *)
    logic[15:0] _e_3678;
    logic[7:0] _e_3682;
    logic[7:0] _e_3683;
    (* src = "src/generated_driver.spade:1140,2" *)
    logic[15:0] _e_3681;
    logic[7:0] _e_3685;
    logic[7:0] _e_3686;
    (* src = "src/generated_driver.spade:1141,2" *)
    logic[15:0] _e_3684;
    logic[7:0] _e_3688;
    logic[7:0] _e_3689;
    (* src = "src/generated_driver.spade:1142,2" *)
    logic[15:0] _e_3687;
    logic[7:0] _e_3691;
    logic[7:0] _e_3692;
    (* src = "src/generated_driver.spade:1143,2" *)
    logic[15:0] _e_3690;
    logic[7:0] _e_3694;
    logic[7:0] _e_3695;
    (* src = "src/generated_driver.spade:1144,2" *)
    logic[15:0] _e_3693;
    logic[7:0] _e_3697;
    logic[7:0] _e_3698;
    (* src = "src/generated_driver.spade:1145,2" *)
    logic[15:0] _e_3696;
    logic[7:0] _e_3700;
    logic[7:0] _e_3701;
    (* src = "src/generated_driver.spade:1146,2" *)
    logic[15:0] _e_3699;
    logic[7:0] _e_3703;
    logic[7:0] _e_3704;
    (* src = "src/generated_driver.spade:1147,2" *)
    logic[15:0] _e_3702;
    logic[7:0] _e_3706;
    logic[7:0] _e_3707;
    (* src = "src/generated_driver.spade:1148,2" *)
    logic[15:0] _e_3705;
    logic[7:0] _e_3709;
    logic[7:0] _e_3710;
    (* src = "src/generated_driver.spade:1149,2" *)
    logic[15:0] _e_3708;
    logic[7:0] _e_3712;
    logic[7:0] _e_3713;
    (* src = "src/generated_driver.spade:1150,2" *)
    logic[15:0] _e_3711;
    logic[7:0] _e_3715;
    logic[7:0] _e_3716;
    (* src = "src/generated_driver.spade:1151,2" *)
    logic[15:0] _e_3714;
    logic[7:0] _e_3718;
    logic[7:0] _e_3719;
    (* src = "src/generated_driver.spade:1152,2" *)
    logic[15:0] _e_3717;
    logic[7:0] _e_3721;
    logic[7:0] _e_3722;
    (* src = "src/generated_driver.spade:1153,2" *)
    logic[15:0] _e_3720;
    logic[7:0] _e_3724;
    logic[7:0] _e_3725;
    (* src = "src/generated_driver.spade:1154,2" *)
    logic[15:0] _e_3723;
    logic[7:0] _e_3727;
    logic[7:0] _e_3728;
    (* src = "src/generated_driver.spade:1155,2" *)
    logic[15:0] _e_3726;
    logic[7:0] _e_3730;
    logic[7:0] _e_3731;
    (* src = "src/generated_driver.spade:1156,2" *)
    logic[15:0] _e_3729;
    logic[7:0] _e_3733;
    logic[7:0] _e_3734;
    (* src = "src/generated_driver.spade:1157,2" *)
    logic[15:0] _e_3732;
    logic[7:0] _e_3736;
    logic[7:0] _e_3737;
    (* src = "src/generated_driver.spade:1158,2" *)
    logic[15:0] _e_3735;
    (* src = "src/generated_driver.spade:34,58" *)
    logic[17999:0] _e_362;
    (* src = "src/generated_driver.spade:34,24" *)
    logic[16-1:0] \commands [1125-1:0];
    (* src = "src/generated_driver.spade:1160,50" *)
    logic[10:0] _e_3741;
    (* src = "src/generated_driver.spade:1160,23" *)
    logic[15:0] \mem_out ;
    logic[7:0] \a ;
    logic[7:0] \b ;
    (* src = "src/generated_driver.spade:1163,9" *)
    logic[15:0] _e_3748;
    always @(posedge \clk ) begin
        \s1_rst  <= \rst ;
    end
    always @(posedge \clk ) begin
        \s1_state  <= \state ;
    end
    always @(posedge \clk ) begin
        \s1_read_idx  <= \read_idx ;
    end
    always @(posedge \clk ) begin
        \s1_mem_out  <= \mem_out ;
    end
    assign _e_307 = 32'd0;
    assign _e_306 = {1'd0, _e_307, 15'bX};
    assign _e_310 = \state [46:15];
    assign _e_3772 = \state [47] == 1'd0;
    assign _e_3774 = 32'd100000000;
    assign _e_3773 = _e_310 == _e_3774;
    assign _e_3775 = _e_3772 && _e_3773;
    assign _e_313 = 0;
    assign _e_314 = 32'd0;
    assign _e_312 = {1'd1, _e_313, _e_314};
    assign \duration  = \state [46:15];
    assign _e_3777 = \state [47] == 1'd0;
    assign _e_3778 = 1;
    assign _e_3779 = _e_3777 && _e_3778;
    assign _e_321 = 32'd1;
    assign _e_319 = $signed(\duration ) + $signed(_e_321);
    assign _e_318 = _e_319[31:0];
    assign _e_317 = {1'd0, _e_318, 15'bX};
    assign _e_322 = \state [46:32];
    assign _e_323 = \state [31:0];
    assign _e_3781 = \state [47] == 1'd1;
    assign _e_3783 = 1124;
    assign _e_3782 = _e_322 == _e_3783;
    assign _e_3785 = 32'd5;
    assign _e_3784 = _e_323 == _e_3785;
    assign _e_3786 = _e_3781 && _e_3782;
    assign _e_3787 = _e_3786 && _e_3784;
    assign _e_327 = 32'd0;
    assign _e_326 = {1'd0, _e_327, 15'bX};
    assign \idx  = \state [46:32];
    assign _e_329 = \state [31:0];
    assign _e_3789 = \state [47] == 1'd1;
    assign _e_3790 = 1;
    assign _e_3792 = 32'd5;
    assign _e_3791 = _e_329 == _e_3792;
    assign _e_3793 = _e_3789 && _e_3790;
    assign _e_3794 = _e_3793 && _e_3791;
    assign _e_336 = 1;
    assign _e_334 = $signed(\idx ) + $signed(_e_336);
    assign _e_333 = _e_334[14:0];
    assign _e_337 = 32'd0;
    assign _e_332 = {1'd1, _e_333, _e_337};
    assign idx_n1 = \state [46:32];
    assign duration_n1 = \state [31:0];
    assign _e_3796 = \state [47] == 1'd1;
    assign _e_3797 = 1;
    assign _e_3798 = 1;
    assign _e_3799 = _e_3796 && _e_3797;
    assign _e_3800 = _e_3799 && _e_3798;
    assign _e_343 = idx_n1[14:0];
    assign _e_348 = 32'd1;
    assign _e_346 = $signed(duration_n1) + $signed(_e_348);
    assign _e_345 = _e_346[31:0];
    assign _e_342 = {1'd1, _e_343, _e_345};
    always_comb begin
        priority casez ({_e_3775, _e_3779, _e_3787, _e_3794, _e_3800})
            5'b1????: _e_308 = _e_312;
            5'b01???: _e_308 = _e_317;
            5'b001??: _e_308 = _e_326;
            5'b0001?: _e_308 = _e_332;
            5'b00001: _e_308 = _e_342;
            5'b?: _e_308 = 'x;
        endcase
    end
    always @(posedge \clk , posedge \rst ) begin
        if (\rst ) begin
            \state  <= _e_306;
        end
        else begin
            \state  <= _e_308;
        end
    end
    assign idx_n2 = \state [46:32];
    assign \_  = \state [31:0];
    assign _e_3802 = \state [47] == 1'd1;
    assign _e_3803 = 1;
    assign _e_3804 = 1;
    assign _e_3805 = _e_3802 && _e_3803;
    assign _e_3806 = _e_3805 && _e_3804;
    assign __n1 = \state [46:15];
    assign _e_3808 = \state [47] == 1'd0;
    assign _e_3809 = 1;
    assign _e_3810 = _e_3808 && _e_3809;
    assign _e_357 = 0;
    always_comb begin
        priority casez ({_e_3806, _e_3810})
            2'b1?: \read_idx  = idx_n2;
            2'b01: \read_idx  = _e_357;
            2'b?: \read_idx  = 'x;
        endcase
    end
    
    assign _e_364 = 0;
    assign _e_365 = 0;
    assign _e_363 = {_e_364, _e_365};
    assign _e_367 = 128;
    assign _e_368 = 0;
    assign _e_366 = {_e_367, _e_368};
    assign _e_370 = 128;
    assign _e_371 = 20;
    assign _e_369 = {_e_370, _e_371};
    assign _e_373 = 128;
    assign _e_374 = 148;
    assign _e_372 = {_e_373, _e_374};
    assign _e_376 = 128;
    assign _e_377 = 20;
    assign _e_375 = {_e_376, _e_377};
    assign _e_379 = 10;
    assign _e_380 = 0;
    assign _e_378 = {_e_379, _e_380};
    assign _e_382 = 138;
    assign _e_383 = 0;
    assign _e_381 = {_e_382, _e_383};
    assign _e_385 = 138;
    assign _e_386 = 50;
    assign _e_384 = {_e_385, _e_386};
    assign _e_388 = 138;
    assign _e_389 = 178;
    assign _e_387 = {_e_388, _e_389};
    assign _e_391 = 138;
    assign _e_392 = 50;
    assign _e_390 = {_e_391, _e_392};
    assign _e_394 = 0;
    assign _e_395 = 0;
    assign _e_393 = {_e_394, _e_395};
    assign _e_397 = 128;
    assign _e_398 = 0;
    assign _e_396 = {_e_397, _e_398};
    assign _e_400 = 128;
    assign _e_401 = 51;
    assign _e_399 = {_e_400, _e_401};
    assign _e_403 = 128;
    assign _e_404 = 179;
    assign _e_402 = {_e_403, _e_404};
    assign _e_406 = 128;
    assign _e_407 = 51;
    assign _e_405 = {_e_406, _e_407};
    assign _e_409 = 20;
    assign _e_410 = 0;
    assign _e_408 = {_e_409, _e_410};
    assign _e_412 = 148;
    assign _e_413 = 0;
    assign _e_411 = {_e_412, _e_413};
    assign _e_415 = 148;
    assign _e_416 = 52;
    assign _e_414 = {_e_415, _e_416};
    assign _e_418 = 148;
    assign _e_419 = 180;
    assign _e_417 = {_e_418, _e_419};
    assign _e_421 = 148;
    assign _e_422 = 52;
    assign _e_420 = {_e_421, _e_422};
    assign _e_424 = 20;
    assign _e_425 = 0;
    assign _e_423 = {_e_424, _e_425};
    assign _e_427 = 148;
    assign _e_428 = 0;
    assign _e_426 = {_e_427, _e_428};
    assign _e_430 = 178;
    assign _e_431 = 61;
    assign _e_429 = {_e_430, _e_431};
    assign _e_433 = 178;
    assign _e_434 = 189;
    assign _e_432 = {_e_433, _e_434};
    assign _e_436 = 178;
    assign _e_437 = 61;
    assign _e_435 = {_e_436, _e_437};
    assign _e_439 = 61;
    assign _e_440 = 0;
    assign _e_438 = {_e_439, _e_440};
    assign _e_442 = 189;
    assign _e_443 = 0;
    assign _e_441 = {_e_442, _e_443};
    assign _e_445 = 189;
    assign _e_446 = 61;
    assign _e_444 = {_e_445, _e_446};
    assign _e_448 = 189;
    assign _e_449 = 189;
    assign _e_447 = {_e_448, _e_449};
    assign _e_451 = 189;
    assign _e_452 = 61;
    assign _e_450 = {_e_451, _e_452};
    assign _e_454 = 61;
    assign _e_455 = 0;
    assign _e_453 = {_e_454, _e_455};
    assign _e_457 = 189;
    assign _e_458 = 0;
    assign _e_456 = {_e_457, _e_458};
    assign _e_460 = 179;
    assign _e_461 = 61;
    assign _e_459 = {_e_460, _e_461};
    assign _e_463 = 179;
    assign _e_464 = 189;
    assign _e_462 = {_e_463, _e_464};
    assign _e_466 = 179;
    assign _e_467 = 61;
    assign _e_465 = {_e_466, _e_467};
    assign _e_469 = 52;
    assign _e_470 = 0;
    assign _e_468 = {_e_469, _e_470};
    assign _e_472 = 180;
    assign _e_473 = 0;
    assign _e_471 = {_e_472, _e_473};
    assign _e_475 = 178;
    assign _e_476 = 62;
    assign _e_474 = {_e_475, _e_476};
    assign _e_478 = 178;
    assign _e_479 = 190;
    assign _e_477 = {_e_478, _e_479};
    assign _e_481 = 178;
    assign _e_482 = 62;
    assign _e_480 = {_e_481, _e_482};
    assign _e_484 = 62;
    assign _e_485 = 0;
    assign _e_483 = {_e_484, _e_485};
    assign _e_487 = 190;
    assign _e_488 = 0;
    assign _e_486 = {_e_487, _e_488};
    assign _e_490 = 190;
    assign _e_491 = 62;
    assign _e_489 = {_e_490, _e_491};
    assign _e_493 = 190;
    assign _e_494 = 190;
    assign _e_492 = {_e_493, _e_494};
    assign _e_496 = 190;
    assign _e_497 = 62;
    assign _e_495 = {_e_496, _e_497};
    assign _e_499 = 62;
    assign _e_500 = 0;
    assign _e_498 = {_e_499, _e_500};
    assign _e_502 = 190;
    assign _e_503 = 0;
    assign _e_501 = {_e_502, _e_503};
    assign _e_505 = 128;
    assign _e_506 = 62;
    assign _e_504 = {_e_505, _e_506};
    assign _e_508 = 128;
    assign _e_509 = 190;
    assign _e_507 = {_e_508, _e_509};
    assign _e_511 = 128;
    assign _e_512 = 62;
    assign _e_510 = {_e_511, _e_512};
    assign _e_514 = 20;
    assign _e_515 = 0;
    assign _e_513 = {_e_514, _e_515};
    assign _e_517 = 148;
    assign _e_518 = 0;
    assign _e_516 = {_e_517, _e_518};
    assign _e_520 = 138;
    assign _e_521 = 63;
    assign _e_519 = {_e_520, _e_521};
    assign _e_523 = 138;
    assign _e_524 = 191;
    assign _e_522 = {_e_523, _e_524};
    assign _e_526 = 138;
    assign _e_527 = 63;
    assign _e_525 = {_e_526, _e_527};
    assign _e_529 = 63;
    assign _e_530 = 0;
    assign _e_528 = {_e_529, _e_530};
    assign _e_532 = 191;
    assign _e_533 = 0;
    assign _e_531 = {_e_532, _e_533};
    assign _e_535 = 191;
    assign _e_536 = 63;
    assign _e_534 = {_e_535, _e_536};
    assign _e_538 = 191;
    assign _e_539 = 191;
    assign _e_537 = {_e_538, _e_539};
    assign _e_541 = 191;
    assign _e_542 = 63;
    assign _e_540 = {_e_541, _e_542};
    assign _e_544 = 63;
    assign _e_545 = 0;
    assign _e_543 = {_e_544, _e_545};
    assign _e_547 = 191;
    assign _e_548 = 0;
    assign _e_546 = {_e_547, _e_548};
    assign _e_550 = 128;
    assign _e_551 = 63;
    assign _e_549 = {_e_550, _e_551};
    assign _e_553 = 128;
    assign _e_554 = 191;
    assign _e_552 = {_e_553, _e_554};
    assign _e_556 = 128;
    assign _e_557 = 63;
    assign _e_555 = {_e_556, _e_557};
    assign _e_559 = 52;
    assign _e_560 = 0;
    assign _e_558 = {_e_559, _e_560};
    assign _e_562 = 180;
    assign _e_563 = 0;
    assign _e_561 = {_e_562, _e_563};
    assign _e_565 = 138;
    assign _e_566 = 64;
    assign _e_564 = {_e_565, _e_566};
    assign _e_568 = 138;
    assign _e_569 = 192;
    assign _e_567 = {_e_568, _e_569};
    assign _e_571 = 138;
    assign _e_572 = 64;
    assign _e_570 = {_e_571, _e_572};
    assign _e_574 = 64;
    assign _e_575 = 0;
    assign _e_573 = {_e_574, _e_575};
    assign _e_577 = 192;
    assign _e_578 = 0;
    assign _e_576 = {_e_577, _e_578};
    assign _e_580 = 192;
    assign _e_581 = 64;
    assign _e_579 = {_e_580, _e_581};
    assign _e_583 = 192;
    assign _e_584 = 192;
    assign _e_582 = {_e_583, _e_584};
    assign _e_586 = 192;
    assign _e_587 = 64;
    assign _e_585 = {_e_586, _e_587};
    assign _e_589 = 64;
    assign _e_590 = 0;
    assign _e_588 = {_e_589, _e_590};
    assign _e_592 = 192;
    assign _e_593 = 0;
    assign _e_591 = {_e_592, _e_593};
    assign _e_595 = 179;
    assign _e_596 = 64;
    assign _e_594 = {_e_595, _e_596};
    assign _e_598 = 179;
    assign _e_599 = 192;
    assign _e_597 = {_e_598, _e_599};
    assign _e_601 = 179;
    assign _e_602 = 64;
    assign _e_600 = {_e_601, _e_602};
    assign _e_604 = 61;
    assign _e_605 = 0;
    assign _e_603 = {_e_604, _e_605};
    assign _e_607 = 189;
    assign _e_608 = 0;
    assign _e_606 = {_e_607, _e_608};
    assign _e_610 = 190;
    assign _e_611 = 127;
    assign _e_609 = {_e_610, _e_611};
    assign _e_613 = 190;
    assign _e_614 = 255;
    assign _e_612 = {_e_613, _e_614};
    assign _e_616 = 190;
    assign _e_617 = 127;
    assign _e_615 = {_e_616, _e_617};
    assign _e_619 = 127;
    assign _e_620 = 0;
    assign _e_618 = {_e_619, _e_620};
    assign _e_622 = 255;
    assign _e_623 = 0;
    assign _e_621 = {_e_622, _e_623};
    assign _e_625 = 255;
    assign _e_626 = 127;
    assign _e_624 = {_e_625, _e_626};
    assign _e_628 = 255;
    assign _e_629 = 255;
    assign _e_627 = {_e_628, _e_629};
    assign _e_631 = 255;
    assign _e_632 = 127;
    assign _e_630 = {_e_631, _e_632};
    assign _e_634 = 63;
    assign _e_635 = 0;
    assign _e_633 = {_e_634, _e_635};
    assign _e_637 = 191;
    assign _e_638 = 0;
    assign _e_636 = {_e_637, _e_638};
    assign _e_640 = 192;
    assign _e_641 = 30;
    assign _e_639 = {_e_640, _e_641};
    assign _e_643 = 192;
    assign _e_644 = 158;
    assign _e_642 = {_e_643, _e_644};
    assign _e_646 = 192;
    assign _e_647 = 30;
    assign _e_645 = {_e_646, _e_647};
    assign _e_649 = 30;
    assign _e_650 = 0;
    assign _e_648 = {_e_649, _e_650};
    assign _e_652 = 158;
    assign _e_653 = 0;
    assign _e_651 = {_e_652, _e_653};
    assign _e_655 = 158;
    assign _e_656 = 30;
    assign _e_654 = {_e_655, _e_656};
    assign _e_658 = 158;
    assign _e_659 = 158;
    assign _e_657 = {_e_658, _e_659};
    assign _e_661 = 158;
    assign _e_662 = 30;
    assign _e_660 = {_e_661, _e_662};
    assign _e_664 = 30;
    assign _e_665 = 0;
    assign _e_663 = {_e_664, _e_665};
    assign _e_667 = 158;
    assign _e_668 = 0;
    assign _e_666 = {_e_667, _e_668};
    assign _e_670 = 255;
    assign _e_671 = 30;
    assign _e_669 = {_e_670, _e_671};
    assign _e_673 = 255;
    assign _e_674 = 158;
    assign _e_672 = {_e_673, _e_674};
    assign _e_676 = 255;
    assign _e_677 = 30;
    assign _e_675 = {_e_676, _e_677};
    assign _e_679 = 10;
    assign _e_680 = 0;
    assign _e_678 = {_e_679, _e_680};
    assign _e_682 = 138;
    assign _e_683 = 0;
    assign _e_681 = {_e_682, _e_683};
    assign _e_685 = 128;
    assign _e_686 = 61;
    assign _e_684 = {_e_685, _e_686};
    assign _e_688 = 128;
    assign _e_689 = 189;
    assign _e_687 = {_e_688, _e_689};
    assign _e_691 = 128;
    assign _e_692 = 61;
    assign _e_690 = {_e_691, _e_692};
    assign _e_694 = 20;
    assign _e_695 = 0;
    assign _e_693 = {_e_694, _e_695};
    assign _e_697 = 148;
    assign _e_698 = 0;
    assign _e_696 = {_e_697, _e_698};
    assign _e_700 = 138;
    assign _e_701 = 62;
    assign _e_699 = {_e_700, _e_701};
    assign _e_703 = 138;
    assign _e_704 = 190;
    assign _e_702 = {_e_703, _e_704};
    assign _e_706 = 138;
    assign _e_707 = 62;
    assign _e_705 = {_e_706, _e_707};
    assign _e_709 = 20;
    assign _e_710 = 0;
    assign _e_708 = {_e_709, _e_710};
    assign _e_712 = 148;
    assign _e_713 = 0;
    assign _e_711 = {_e_712, _e_713};
    assign _e_715 = 128;
    assign _e_716 = 63;
    assign _e_714 = {_e_715, _e_716};
    assign _e_718 = 128;
    assign _e_719 = 191;
    assign _e_717 = {_e_718, _e_719};
    assign _e_721 = 128;
    assign _e_722 = 63;
    assign _e_720 = {_e_721, _e_722};
    assign _e_724 = 61;
    assign _e_725 = 0;
    assign _e_723 = {_e_724, _e_725};
    assign _e_727 = 189;
    assign _e_728 = 0;
    assign _e_726 = {_e_727, _e_728};
    assign _e_730 = 190;
    assign _e_731 = 20;
    assign _e_729 = {_e_730, _e_731};
    assign _e_733 = 190;
    assign _e_734 = 148;
    assign _e_732 = {_e_733, _e_734};
    assign _e_736 = 190;
    assign _e_737 = 20;
    assign _e_735 = {_e_736, _e_737};
    assign _e_739 = 20;
    assign _e_740 = 0;
    assign _e_738 = {_e_739, _e_740};
    assign _e_742 = 148;
    assign _e_743 = 0;
    assign _e_741 = {_e_742, _e_743};
    assign _e_745 = 148;
    assign _e_746 = 20;
    assign _e_744 = {_e_745, _e_746};
    assign _e_748 = 148;
    assign _e_749 = 148;
    assign _e_747 = {_e_748, _e_749};
    assign _e_751 = 148;
    assign _e_752 = 20;
    assign _e_750 = {_e_751, _e_752};
    assign _e_754 = 20;
    assign _e_755 = 0;
    assign _e_753 = {_e_754, _e_755};
    assign _e_757 = 148;
    assign _e_758 = 0;
    assign _e_756 = {_e_757, _e_758};
    assign _e_760 = 191;
    assign _e_761 = 20;
    assign _e_759 = {_e_760, _e_761};
    assign _e_763 = 191;
    assign _e_764 = 148;
    assign _e_762 = {_e_763, _e_764};
    assign _e_766 = 191;
    assign _e_767 = 20;
    assign _e_765 = {_e_766, _e_767};
    assign _e_769 = 11;
    assign _e_770 = 0;
    assign _e_768 = {_e_769, _e_770};
    assign _e_772 = 139;
    assign _e_773 = 0;
    assign _e_771 = {_e_772, _e_773};
    assign _e_775 = 139;
    assign _e_776 = 50;
    assign _e_774 = {_e_775, _e_776};
    assign _e_778 = 139;
    assign _e_779 = 178;
    assign _e_777 = {_e_778, _e_779};
    assign _e_781 = 139;
    assign _e_782 = 50;
    assign _e_780 = {_e_781, _e_782};
    assign _e_784 = 0;
    assign _e_785 = 0;
    assign _e_783 = {_e_784, _e_785};
    assign _e_787 = 128;
    assign _e_788 = 0;
    assign _e_786 = {_e_787, _e_788};
    assign _e_790 = 128;
    assign _e_791 = 51;
    assign _e_789 = {_e_790, _e_791};
    assign _e_793 = 128;
    assign _e_794 = 179;
    assign _e_792 = {_e_793, _e_794};
    assign _e_796 = 128;
    assign _e_797 = 51;
    assign _e_795 = {_e_796, _e_797};
    assign _e_799 = 20;
    assign _e_800 = 0;
    assign _e_798 = {_e_799, _e_800};
    assign _e_802 = 148;
    assign _e_803 = 0;
    assign _e_801 = {_e_802, _e_803};
    assign _e_805 = 148;
    assign _e_806 = 52;
    assign _e_804 = {_e_805, _e_806};
    assign _e_808 = 148;
    assign _e_809 = 180;
    assign _e_807 = {_e_808, _e_809};
    assign _e_811 = 148;
    assign _e_812 = 52;
    assign _e_810 = {_e_811, _e_812};
    assign _e_814 = 20;
    assign _e_815 = 0;
    assign _e_813 = {_e_814, _e_815};
    assign _e_817 = 148;
    assign _e_818 = 0;
    assign _e_816 = {_e_817, _e_818};
    assign _e_820 = 178;
    assign _e_821 = 61;
    assign _e_819 = {_e_820, _e_821};
    assign _e_823 = 178;
    assign _e_824 = 189;
    assign _e_822 = {_e_823, _e_824};
    assign _e_826 = 178;
    assign _e_827 = 61;
    assign _e_825 = {_e_826, _e_827};
    assign _e_829 = 61;
    assign _e_830 = 0;
    assign _e_828 = {_e_829, _e_830};
    assign _e_832 = 189;
    assign _e_833 = 0;
    assign _e_831 = {_e_832, _e_833};
    assign _e_835 = 189;
    assign _e_836 = 61;
    assign _e_834 = {_e_835, _e_836};
    assign _e_838 = 189;
    assign _e_839 = 189;
    assign _e_837 = {_e_838, _e_839};
    assign _e_841 = 189;
    assign _e_842 = 61;
    assign _e_840 = {_e_841, _e_842};
    assign _e_844 = 61;
    assign _e_845 = 0;
    assign _e_843 = {_e_844, _e_845};
    assign _e_847 = 189;
    assign _e_848 = 0;
    assign _e_846 = {_e_847, _e_848};
    assign _e_850 = 179;
    assign _e_851 = 61;
    assign _e_849 = {_e_850, _e_851};
    assign _e_853 = 179;
    assign _e_854 = 189;
    assign _e_852 = {_e_853, _e_854};
    assign _e_856 = 179;
    assign _e_857 = 61;
    assign _e_855 = {_e_856, _e_857};
    assign _e_859 = 52;
    assign _e_860 = 0;
    assign _e_858 = {_e_859, _e_860};
    assign _e_862 = 180;
    assign _e_863 = 0;
    assign _e_861 = {_e_862, _e_863};
    assign _e_865 = 178;
    assign _e_866 = 62;
    assign _e_864 = {_e_865, _e_866};
    assign _e_868 = 178;
    assign _e_869 = 190;
    assign _e_867 = {_e_868, _e_869};
    assign _e_871 = 178;
    assign _e_872 = 62;
    assign _e_870 = {_e_871, _e_872};
    assign _e_874 = 62;
    assign _e_875 = 0;
    assign _e_873 = {_e_874, _e_875};
    assign _e_877 = 190;
    assign _e_878 = 0;
    assign _e_876 = {_e_877, _e_878};
    assign _e_880 = 190;
    assign _e_881 = 62;
    assign _e_879 = {_e_880, _e_881};
    assign _e_883 = 190;
    assign _e_884 = 190;
    assign _e_882 = {_e_883, _e_884};
    assign _e_886 = 190;
    assign _e_887 = 62;
    assign _e_885 = {_e_886, _e_887};
    assign _e_889 = 62;
    assign _e_890 = 0;
    assign _e_888 = {_e_889, _e_890};
    assign _e_892 = 190;
    assign _e_893 = 0;
    assign _e_891 = {_e_892, _e_893};
    assign _e_895 = 128;
    assign _e_896 = 62;
    assign _e_894 = {_e_895, _e_896};
    assign _e_898 = 128;
    assign _e_899 = 190;
    assign _e_897 = {_e_898, _e_899};
    assign _e_901 = 128;
    assign _e_902 = 62;
    assign _e_900 = {_e_901, _e_902};
    assign _e_904 = 20;
    assign _e_905 = 0;
    assign _e_903 = {_e_904, _e_905};
    assign _e_907 = 148;
    assign _e_908 = 0;
    assign _e_906 = {_e_907, _e_908};
    assign _e_910 = 139;
    assign _e_911 = 63;
    assign _e_909 = {_e_910, _e_911};
    assign _e_913 = 139;
    assign _e_914 = 191;
    assign _e_912 = {_e_913, _e_914};
    assign _e_916 = 139;
    assign _e_917 = 63;
    assign _e_915 = {_e_916, _e_917};
    assign _e_919 = 63;
    assign _e_920 = 0;
    assign _e_918 = {_e_919, _e_920};
    assign _e_922 = 191;
    assign _e_923 = 0;
    assign _e_921 = {_e_922, _e_923};
    assign _e_925 = 191;
    assign _e_926 = 63;
    assign _e_924 = {_e_925, _e_926};
    assign _e_928 = 191;
    assign _e_929 = 191;
    assign _e_927 = {_e_928, _e_929};
    assign _e_931 = 191;
    assign _e_932 = 63;
    assign _e_930 = {_e_931, _e_932};
    assign _e_934 = 63;
    assign _e_935 = 0;
    assign _e_933 = {_e_934, _e_935};
    assign _e_937 = 191;
    assign _e_938 = 0;
    assign _e_936 = {_e_937, _e_938};
    assign _e_940 = 128;
    assign _e_941 = 63;
    assign _e_939 = {_e_940, _e_941};
    assign _e_943 = 128;
    assign _e_944 = 191;
    assign _e_942 = {_e_943, _e_944};
    assign _e_946 = 128;
    assign _e_947 = 63;
    assign _e_945 = {_e_946, _e_947};
    assign _e_949 = 52;
    assign _e_950 = 0;
    assign _e_948 = {_e_949, _e_950};
    assign _e_952 = 180;
    assign _e_953 = 0;
    assign _e_951 = {_e_952, _e_953};
    assign _e_955 = 139;
    assign _e_956 = 64;
    assign _e_954 = {_e_955, _e_956};
    assign _e_958 = 139;
    assign _e_959 = 192;
    assign _e_957 = {_e_958, _e_959};
    assign _e_961 = 139;
    assign _e_962 = 64;
    assign _e_960 = {_e_961, _e_962};
    assign _e_964 = 64;
    assign _e_965 = 0;
    assign _e_963 = {_e_964, _e_965};
    assign _e_967 = 192;
    assign _e_968 = 0;
    assign _e_966 = {_e_967, _e_968};
    assign _e_970 = 192;
    assign _e_971 = 64;
    assign _e_969 = {_e_970, _e_971};
    assign _e_973 = 192;
    assign _e_974 = 192;
    assign _e_972 = {_e_973, _e_974};
    assign _e_976 = 192;
    assign _e_977 = 64;
    assign _e_975 = {_e_976, _e_977};
    assign _e_979 = 64;
    assign _e_980 = 0;
    assign _e_978 = {_e_979, _e_980};
    assign _e_982 = 192;
    assign _e_983 = 0;
    assign _e_981 = {_e_982, _e_983};
    assign _e_985 = 179;
    assign _e_986 = 64;
    assign _e_984 = {_e_985, _e_986};
    assign _e_988 = 179;
    assign _e_989 = 192;
    assign _e_987 = {_e_988, _e_989};
    assign _e_991 = 179;
    assign _e_992 = 64;
    assign _e_990 = {_e_991, _e_992};
    assign _e_994 = 61;
    assign _e_995 = 0;
    assign _e_993 = {_e_994, _e_995};
    assign _e_997 = 189;
    assign _e_998 = 0;
    assign _e_996 = {_e_997, _e_998};
    assign _e_1000 = 190;
    assign _e_1001 = 127;
    assign _e_999 = {_e_1000, _e_1001};
    assign _e_1003 = 190;
    assign _e_1004 = 255;
    assign _e_1002 = {_e_1003, _e_1004};
    assign _e_1006 = 190;
    assign _e_1007 = 127;
    assign _e_1005 = {_e_1006, _e_1007};
    assign _e_1009 = 127;
    assign _e_1010 = 0;
    assign _e_1008 = {_e_1009, _e_1010};
    assign _e_1012 = 255;
    assign _e_1013 = 0;
    assign _e_1011 = {_e_1012, _e_1013};
    assign _e_1015 = 255;
    assign _e_1016 = 127;
    assign _e_1014 = {_e_1015, _e_1016};
    assign _e_1018 = 255;
    assign _e_1019 = 255;
    assign _e_1017 = {_e_1018, _e_1019};
    assign _e_1021 = 255;
    assign _e_1022 = 127;
    assign _e_1020 = {_e_1021, _e_1022};
    assign _e_1024 = 63;
    assign _e_1025 = 0;
    assign _e_1023 = {_e_1024, _e_1025};
    assign _e_1027 = 191;
    assign _e_1028 = 0;
    assign _e_1026 = {_e_1027, _e_1028};
    assign _e_1030 = 192;
    assign _e_1031 = 31;
    assign _e_1029 = {_e_1030, _e_1031};
    assign _e_1033 = 192;
    assign _e_1034 = 159;
    assign _e_1032 = {_e_1033, _e_1034};
    assign _e_1036 = 192;
    assign _e_1037 = 31;
    assign _e_1035 = {_e_1036, _e_1037};
    assign _e_1039 = 31;
    assign _e_1040 = 0;
    assign _e_1038 = {_e_1039, _e_1040};
    assign _e_1042 = 159;
    assign _e_1043 = 0;
    assign _e_1041 = {_e_1042, _e_1043};
    assign _e_1045 = 159;
    assign _e_1046 = 31;
    assign _e_1044 = {_e_1045, _e_1046};
    assign _e_1048 = 159;
    assign _e_1049 = 159;
    assign _e_1047 = {_e_1048, _e_1049};
    assign _e_1051 = 159;
    assign _e_1052 = 31;
    assign _e_1050 = {_e_1051, _e_1052};
    assign _e_1054 = 31;
    assign _e_1055 = 0;
    assign _e_1053 = {_e_1054, _e_1055};
    assign _e_1057 = 159;
    assign _e_1058 = 0;
    assign _e_1056 = {_e_1057, _e_1058};
    assign _e_1060 = 255;
    assign _e_1061 = 31;
    assign _e_1059 = {_e_1060, _e_1061};
    assign _e_1063 = 255;
    assign _e_1064 = 159;
    assign _e_1062 = {_e_1063, _e_1064};
    assign _e_1066 = 255;
    assign _e_1067 = 31;
    assign _e_1065 = {_e_1066, _e_1067};
    assign _e_1069 = 11;
    assign _e_1070 = 0;
    assign _e_1068 = {_e_1069, _e_1070};
    assign _e_1072 = 139;
    assign _e_1073 = 0;
    assign _e_1071 = {_e_1072, _e_1073};
    assign _e_1075 = 128;
    assign _e_1076 = 61;
    assign _e_1074 = {_e_1075, _e_1076};
    assign _e_1078 = 128;
    assign _e_1079 = 189;
    assign _e_1077 = {_e_1078, _e_1079};
    assign _e_1081 = 128;
    assign _e_1082 = 61;
    assign _e_1080 = {_e_1081, _e_1082};
    assign _e_1084 = 20;
    assign _e_1085 = 0;
    assign _e_1083 = {_e_1084, _e_1085};
    assign _e_1087 = 148;
    assign _e_1088 = 0;
    assign _e_1086 = {_e_1087, _e_1088};
    assign _e_1090 = 139;
    assign _e_1091 = 62;
    assign _e_1089 = {_e_1090, _e_1091};
    assign _e_1093 = 139;
    assign _e_1094 = 190;
    assign _e_1092 = {_e_1093, _e_1094};
    assign _e_1096 = 139;
    assign _e_1097 = 62;
    assign _e_1095 = {_e_1096, _e_1097};
    assign _e_1099 = 20;
    assign _e_1100 = 0;
    assign _e_1098 = {_e_1099, _e_1100};
    assign _e_1102 = 148;
    assign _e_1103 = 0;
    assign _e_1101 = {_e_1102, _e_1103};
    assign _e_1105 = 128;
    assign _e_1106 = 63;
    assign _e_1104 = {_e_1105, _e_1106};
    assign _e_1108 = 128;
    assign _e_1109 = 191;
    assign _e_1107 = {_e_1108, _e_1109};
    assign _e_1111 = 128;
    assign _e_1112 = 63;
    assign _e_1110 = {_e_1111, _e_1112};
    assign _e_1114 = 61;
    assign _e_1115 = 0;
    assign _e_1113 = {_e_1114, _e_1115};
    assign _e_1117 = 189;
    assign _e_1118 = 0;
    assign _e_1116 = {_e_1117, _e_1118};
    assign _e_1120 = 190;
    assign _e_1121 = 20;
    assign _e_1119 = {_e_1120, _e_1121};
    assign _e_1123 = 190;
    assign _e_1124 = 148;
    assign _e_1122 = {_e_1123, _e_1124};
    assign _e_1126 = 190;
    assign _e_1127 = 20;
    assign _e_1125 = {_e_1126, _e_1127};
    assign _e_1129 = 20;
    assign _e_1130 = 0;
    assign _e_1128 = {_e_1129, _e_1130};
    assign _e_1132 = 148;
    assign _e_1133 = 0;
    assign _e_1131 = {_e_1132, _e_1133};
    assign _e_1135 = 148;
    assign _e_1136 = 20;
    assign _e_1134 = {_e_1135, _e_1136};
    assign _e_1138 = 148;
    assign _e_1139 = 148;
    assign _e_1137 = {_e_1138, _e_1139};
    assign _e_1141 = 148;
    assign _e_1142 = 20;
    assign _e_1140 = {_e_1141, _e_1142};
    assign _e_1144 = 20;
    assign _e_1145 = 0;
    assign _e_1143 = {_e_1144, _e_1145};
    assign _e_1147 = 148;
    assign _e_1148 = 0;
    assign _e_1146 = {_e_1147, _e_1148};
    assign _e_1150 = 191;
    assign _e_1151 = 20;
    assign _e_1149 = {_e_1150, _e_1151};
    assign _e_1153 = 191;
    assign _e_1154 = 148;
    assign _e_1152 = {_e_1153, _e_1154};
    assign _e_1156 = 191;
    assign _e_1157 = 20;
    assign _e_1155 = {_e_1156, _e_1157};
    assign _e_1159 = 12;
    assign _e_1160 = 0;
    assign _e_1158 = {_e_1159, _e_1160};
    assign _e_1162 = 140;
    assign _e_1163 = 0;
    assign _e_1161 = {_e_1162, _e_1163};
    assign _e_1165 = 140;
    assign _e_1166 = 50;
    assign _e_1164 = {_e_1165, _e_1166};
    assign _e_1168 = 140;
    assign _e_1169 = 178;
    assign _e_1167 = {_e_1168, _e_1169};
    assign _e_1171 = 140;
    assign _e_1172 = 50;
    assign _e_1170 = {_e_1171, _e_1172};
    assign _e_1174 = 0;
    assign _e_1175 = 0;
    assign _e_1173 = {_e_1174, _e_1175};
    assign _e_1177 = 128;
    assign _e_1178 = 0;
    assign _e_1176 = {_e_1177, _e_1178};
    assign _e_1180 = 128;
    assign _e_1181 = 51;
    assign _e_1179 = {_e_1180, _e_1181};
    assign _e_1183 = 128;
    assign _e_1184 = 179;
    assign _e_1182 = {_e_1183, _e_1184};
    assign _e_1186 = 128;
    assign _e_1187 = 51;
    assign _e_1185 = {_e_1186, _e_1187};
    assign _e_1189 = 20;
    assign _e_1190 = 0;
    assign _e_1188 = {_e_1189, _e_1190};
    assign _e_1192 = 148;
    assign _e_1193 = 0;
    assign _e_1191 = {_e_1192, _e_1193};
    assign _e_1195 = 148;
    assign _e_1196 = 52;
    assign _e_1194 = {_e_1195, _e_1196};
    assign _e_1198 = 148;
    assign _e_1199 = 180;
    assign _e_1197 = {_e_1198, _e_1199};
    assign _e_1201 = 148;
    assign _e_1202 = 52;
    assign _e_1200 = {_e_1201, _e_1202};
    assign _e_1204 = 20;
    assign _e_1205 = 0;
    assign _e_1203 = {_e_1204, _e_1205};
    assign _e_1207 = 148;
    assign _e_1208 = 0;
    assign _e_1206 = {_e_1207, _e_1208};
    assign _e_1210 = 178;
    assign _e_1211 = 61;
    assign _e_1209 = {_e_1210, _e_1211};
    assign _e_1213 = 178;
    assign _e_1214 = 189;
    assign _e_1212 = {_e_1213, _e_1214};
    assign _e_1216 = 178;
    assign _e_1217 = 61;
    assign _e_1215 = {_e_1216, _e_1217};
    assign _e_1219 = 61;
    assign _e_1220 = 0;
    assign _e_1218 = {_e_1219, _e_1220};
    assign _e_1222 = 189;
    assign _e_1223 = 0;
    assign _e_1221 = {_e_1222, _e_1223};
    assign _e_1225 = 189;
    assign _e_1226 = 61;
    assign _e_1224 = {_e_1225, _e_1226};
    assign _e_1228 = 189;
    assign _e_1229 = 189;
    assign _e_1227 = {_e_1228, _e_1229};
    assign _e_1231 = 189;
    assign _e_1232 = 61;
    assign _e_1230 = {_e_1231, _e_1232};
    assign _e_1234 = 61;
    assign _e_1235 = 0;
    assign _e_1233 = {_e_1234, _e_1235};
    assign _e_1237 = 189;
    assign _e_1238 = 0;
    assign _e_1236 = {_e_1237, _e_1238};
    assign _e_1240 = 179;
    assign _e_1241 = 61;
    assign _e_1239 = {_e_1240, _e_1241};
    assign _e_1243 = 179;
    assign _e_1244 = 189;
    assign _e_1242 = {_e_1243, _e_1244};
    assign _e_1246 = 179;
    assign _e_1247 = 61;
    assign _e_1245 = {_e_1246, _e_1247};
    assign _e_1249 = 52;
    assign _e_1250 = 0;
    assign _e_1248 = {_e_1249, _e_1250};
    assign _e_1252 = 180;
    assign _e_1253 = 0;
    assign _e_1251 = {_e_1252, _e_1253};
    assign _e_1255 = 178;
    assign _e_1256 = 62;
    assign _e_1254 = {_e_1255, _e_1256};
    assign _e_1258 = 178;
    assign _e_1259 = 190;
    assign _e_1257 = {_e_1258, _e_1259};
    assign _e_1261 = 178;
    assign _e_1262 = 62;
    assign _e_1260 = {_e_1261, _e_1262};
    assign _e_1264 = 62;
    assign _e_1265 = 0;
    assign _e_1263 = {_e_1264, _e_1265};
    assign _e_1267 = 190;
    assign _e_1268 = 0;
    assign _e_1266 = {_e_1267, _e_1268};
    assign _e_1270 = 190;
    assign _e_1271 = 62;
    assign _e_1269 = {_e_1270, _e_1271};
    assign _e_1273 = 190;
    assign _e_1274 = 190;
    assign _e_1272 = {_e_1273, _e_1274};
    assign _e_1276 = 190;
    assign _e_1277 = 62;
    assign _e_1275 = {_e_1276, _e_1277};
    assign _e_1279 = 62;
    assign _e_1280 = 0;
    assign _e_1278 = {_e_1279, _e_1280};
    assign _e_1282 = 190;
    assign _e_1283 = 0;
    assign _e_1281 = {_e_1282, _e_1283};
    assign _e_1285 = 128;
    assign _e_1286 = 62;
    assign _e_1284 = {_e_1285, _e_1286};
    assign _e_1288 = 128;
    assign _e_1289 = 190;
    assign _e_1287 = {_e_1288, _e_1289};
    assign _e_1291 = 128;
    assign _e_1292 = 62;
    assign _e_1290 = {_e_1291, _e_1292};
    assign _e_1294 = 20;
    assign _e_1295 = 0;
    assign _e_1293 = {_e_1294, _e_1295};
    assign _e_1297 = 148;
    assign _e_1298 = 0;
    assign _e_1296 = {_e_1297, _e_1298};
    assign _e_1300 = 140;
    assign _e_1301 = 63;
    assign _e_1299 = {_e_1300, _e_1301};
    assign _e_1303 = 140;
    assign _e_1304 = 191;
    assign _e_1302 = {_e_1303, _e_1304};
    assign _e_1306 = 140;
    assign _e_1307 = 63;
    assign _e_1305 = {_e_1306, _e_1307};
    assign _e_1309 = 63;
    assign _e_1310 = 0;
    assign _e_1308 = {_e_1309, _e_1310};
    assign _e_1312 = 191;
    assign _e_1313 = 0;
    assign _e_1311 = {_e_1312, _e_1313};
    assign _e_1315 = 191;
    assign _e_1316 = 63;
    assign _e_1314 = {_e_1315, _e_1316};
    assign _e_1318 = 191;
    assign _e_1319 = 191;
    assign _e_1317 = {_e_1318, _e_1319};
    assign _e_1321 = 191;
    assign _e_1322 = 63;
    assign _e_1320 = {_e_1321, _e_1322};
    assign _e_1324 = 63;
    assign _e_1325 = 0;
    assign _e_1323 = {_e_1324, _e_1325};
    assign _e_1327 = 191;
    assign _e_1328 = 0;
    assign _e_1326 = {_e_1327, _e_1328};
    assign _e_1330 = 128;
    assign _e_1331 = 63;
    assign _e_1329 = {_e_1330, _e_1331};
    assign _e_1333 = 128;
    assign _e_1334 = 191;
    assign _e_1332 = {_e_1333, _e_1334};
    assign _e_1336 = 128;
    assign _e_1337 = 63;
    assign _e_1335 = {_e_1336, _e_1337};
    assign _e_1339 = 52;
    assign _e_1340 = 0;
    assign _e_1338 = {_e_1339, _e_1340};
    assign _e_1342 = 180;
    assign _e_1343 = 0;
    assign _e_1341 = {_e_1342, _e_1343};
    assign _e_1345 = 140;
    assign _e_1346 = 64;
    assign _e_1344 = {_e_1345, _e_1346};
    assign _e_1348 = 140;
    assign _e_1349 = 192;
    assign _e_1347 = {_e_1348, _e_1349};
    assign _e_1351 = 140;
    assign _e_1352 = 64;
    assign _e_1350 = {_e_1351, _e_1352};
    assign _e_1354 = 64;
    assign _e_1355 = 0;
    assign _e_1353 = {_e_1354, _e_1355};
    assign _e_1357 = 192;
    assign _e_1358 = 0;
    assign _e_1356 = {_e_1357, _e_1358};
    assign _e_1360 = 192;
    assign _e_1361 = 64;
    assign _e_1359 = {_e_1360, _e_1361};
    assign _e_1363 = 192;
    assign _e_1364 = 192;
    assign _e_1362 = {_e_1363, _e_1364};
    assign _e_1366 = 192;
    assign _e_1367 = 64;
    assign _e_1365 = {_e_1366, _e_1367};
    assign _e_1369 = 64;
    assign _e_1370 = 0;
    assign _e_1368 = {_e_1369, _e_1370};
    assign _e_1372 = 192;
    assign _e_1373 = 0;
    assign _e_1371 = {_e_1372, _e_1373};
    assign _e_1375 = 179;
    assign _e_1376 = 64;
    assign _e_1374 = {_e_1375, _e_1376};
    assign _e_1378 = 179;
    assign _e_1379 = 192;
    assign _e_1377 = {_e_1378, _e_1379};
    assign _e_1381 = 179;
    assign _e_1382 = 64;
    assign _e_1380 = {_e_1381, _e_1382};
    assign _e_1384 = 61;
    assign _e_1385 = 0;
    assign _e_1383 = {_e_1384, _e_1385};
    assign _e_1387 = 189;
    assign _e_1388 = 0;
    assign _e_1386 = {_e_1387, _e_1388};
    assign _e_1390 = 190;
    assign _e_1391 = 127;
    assign _e_1389 = {_e_1390, _e_1391};
    assign _e_1393 = 190;
    assign _e_1394 = 255;
    assign _e_1392 = {_e_1393, _e_1394};
    assign _e_1396 = 190;
    assign _e_1397 = 127;
    assign _e_1395 = {_e_1396, _e_1397};
    assign _e_1399 = 127;
    assign _e_1400 = 0;
    assign _e_1398 = {_e_1399, _e_1400};
    assign _e_1402 = 255;
    assign _e_1403 = 0;
    assign _e_1401 = {_e_1402, _e_1403};
    assign _e_1405 = 255;
    assign _e_1406 = 127;
    assign _e_1404 = {_e_1405, _e_1406};
    assign _e_1408 = 255;
    assign _e_1409 = 255;
    assign _e_1407 = {_e_1408, _e_1409};
    assign _e_1411 = 255;
    assign _e_1412 = 127;
    assign _e_1410 = {_e_1411, _e_1412};
    assign _e_1414 = 63;
    assign _e_1415 = 0;
    assign _e_1413 = {_e_1414, _e_1415};
    assign _e_1417 = 191;
    assign _e_1418 = 0;
    assign _e_1416 = {_e_1417, _e_1418};
    assign _e_1420 = 192;
    assign _e_1421 = 32;
    assign _e_1419 = {_e_1420, _e_1421};
    assign _e_1423 = 192;
    assign _e_1424 = 160;
    assign _e_1422 = {_e_1423, _e_1424};
    assign _e_1426 = 192;
    assign _e_1427 = 32;
    assign _e_1425 = {_e_1426, _e_1427};
    assign _e_1429 = 32;
    assign _e_1430 = 0;
    assign _e_1428 = {_e_1429, _e_1430};
    assign _e_1432 = 160;
    assign _e_1433 = 0;
    assign _e_1431 = {_e_1432, _e_1433};
    assign _e_1435 = 160;
    assign _e_1436 = 32;
    assign _e_1434 = {_e_1435, _e_1436};
    assign _e_1438 = 160;
    assign _e_1439 = 160;
    assign _e_1437 = {_e_1438, _e_1439};
    assign _e_1441 = 160;
    assign _e_1442 = 32;
    assign _e_1440 = {_e_1441, _e_1442};
    assign _e_1444 = 32;
    assign _e_1445 = 0;
    assign _e_1443 = {_e_1444, _e_1445};
    assign _e_1447 = 160;
    assign _e_1448 = 0;
    assign _e_1446 = {_e_1447, _e_1448};
    assign _e_1450 = 255;
    assign _e_1451 = 32;
    assign _e_1449 = {_e_1450, _e_1451};
    assign _e_1453 = 255;
    assign _e_1454 = 160;
    assign _e_1452 = {_e_1453, _e_1454};
    assign _e_1456 = 255;
    assign _e_1457 = 32;
    assign _e_1455 = {_e_1456, _e_1457};
    assign _e_1459 = 12;
    assign _e_1460 = 0;
    assign _e_1458 = {_e_1459, _e_1460};
    assign _e_1462 = 140;
    assign _e_1463 = 0;
    assign _e_1461 = {_e_1462, _e_1463};
    assign _e_1465 = 128;
    assign _e_1466 = 61;
    assign _e_1464 = {_e_1465, _e_1466};
    assign _e_1468 = 128;
    assign _e_1469 = 189;
    assign _e_1467 = {_e_1468, _e_1469};
    assign _e_1471 = 128;
    assign _e_1472 = 61;
    assign _e_1470 = {_e_1471, _e_1472};
    assign _e_1474 = 20;
    assign _e_1475 = 0;
    assign _e_1473 = {_e_1474, _e_1475};
    assign _e_1477 = 148;
    assign _e_1478 = 0;
    assign _e_1476 = {_e_1477, _e_1478};
    assign _e_1480 = 140;
    assign _e_1481 = 62;
    assign _e_1479 = {_e_1480, _e_1481};
    assign _e_1483 = 140;
    assign _e_1484 = 190;
    assign _e_1482 = {_e_1483, _e_1484};
    assign _e_1486 = 140;
    assign _e_1487 = 62;
    assign _e_1485 = {_e_1486, _e_1487};
    assign _e_1489 = 20;
    assign _e_1490 = 0;
    assign _e_1488 = {_e_1489, _e_1490};
    assign _e_1492 = 148;
    assign _e_1493 = 0;
    assign _e_1491 = {_e_1492, _e_1493};
    assign _e_1495 = 128;
    assign _e_1496 = 63;
    assign _e_1494 = {_e_1495, _e_1496};
    assign _e_1498 = 128;
    assign _e_1499 = 191;
    assign _e_1497 = {_e_1498, _e_1499};
    assign _e_1501 = 128;
    assign _e_1502 = 63;
    assign _e_1500 = {_e_1501, _e_1502};
    assign _e_1504 = 61;
    assign _e_1505 = 0;
    assign _e_1503 = {_e_1504, _e_1505};
    assign _e_1507 = 189;
    assign _e_1508 = 0;
    assign _e_1506 = {_e_1507, _e_1508};
    assign _e_1510 = 190;
    assign _e_1511 = 20;
    assign _e_1509 = {_e_1510, _e_1511};
    assign _e_1513 = 190;
    assign _e_1514 = 148;
    assign _e_1512 = {_e_1513, _e_1514};
    assign _e_1516 = 190;
    assign _e_1517 = 20;
    assign _e_1515 = {_e_1516, _e_1517};
    assign _e_1519 = 20;
    assign _e_1520 = 0;
    assign _e_1518 = {_e_1519, _e_1520};
    assign _e_1522 = 148;
    assign _e_1523 = 0;
    assign _e_1521 = {_e_1522, _e_1523};
    assign _e_1525 = 148;
    assign _e_1526 = 20;
    assign _e_1524 = {_e_1525, _e_1526};
    assign _e_1528 = 148;
    assign _e_1529 = 148;
    assign _e_1527 = {_e_1528, _e_1529};
    assign _e_1531 = 148;
    assign _e_1532 = 20;
    assign _e_1530 = {_e_1531, _e_1532};
    assign _e_1534 = 20;
    assign _e_1535 = 0;
    assign _e_1533 = {_e_1534, _e_1535};
    assign _e_1537 = 148;
    assign _e_1538 = 0;
    assign _e_1536 = {_e_1537, _e_1538};
    assign _e_1540 = 191;
    assign _e_1541 = 20;
    assign _e_1539 = {_e_1540, _e_1541};
    assign _e_1543 = 191;
    assign _e_1544 = 148;
    assign _e_1542 = {_e_1543, _e_1544};
    assign _e_1546 = 191;
    assign _e_1547 = 20;
    assign _e_1545 = {_e_1546, _e_1547};
    assign _e_1549 = 13;
    assign _e_1550 = 0;
    assign _e_1548 = {_e_1549, _e_1550};
    assign _e_1552 = 141;
    assign _e_1553 = 0;
    assign _e_1551 = {_e_1552, _e_1553};
    assign _e_1555 = 141;
    assign _e_1556 = 50;
    assign _e_1554 = {_e_1555, _e_1556};
    assign _e_1558 = 141;
    assign _e_1559 = 178;
    assign _e_1557 = {_e_1558, _e_1559};
    assign _e_1561 = 141;
    assign _e_1562 = 50;
    assign _e_1560 = {_e_1561, _e_1562};
    assign _e_1564 = 0;
    assign _e_1565 = 0;
    assign _e_1563 = {_e_1564, _e_1565};
    assign _e_1567 = 128;
    assign _e_1568 = 0;
    assign _e_1566 = {_e_1567, _e_1568};
    assign _e_1570 = 128;
    assign _e_1571 = 51;
    assign _e_1569 = {_e_1570, _e_1571};
    assign _e_1573 = 128;
    assign _e_1574 = 179;
    assign _e_1572 = {_e_1573, _e_1574};
    assign _e_1576 = 128;
    assign _e_1577 = 51;
    assign _e_1575 = {_e_1576, _e_1577};
    assign _e_1579 = 20;
    assign _e_1580 = 0;
    assign _e_1578 = {_e_1579, _e_1580};
    assign _e_1582 = 148;
    assign _e_1583 = 0;
    assign _e_1581 = {_e_1582, _e_1583};
    assign _e_1585 = 148;
    assign _e_1586 = 52;
    assign _e_1584 = {_e_1585, _e_1586};
    assign _e_1588 = 148;
    assign _e_1589 = 180;
    assign _e_1587 = {_e_1588, _e_1589};
    assign _e_1591 = 148;
    assign _e_1592 = 52;
    assign _e_1590 = {_e_1591, _e_1592};
    assign _e_1594 = 20;
    assign _e_1595 = 0;
    assign _e_1593 = {_e_1594, _e_1595};
    assign _e_1597 = 148;
    assign _e_1598 = 0;
    assign _e_1596 = {_e_1597, _e_1598};
    assign _e_1600 = 178;
    assign _e_1601 = 61;
    assign _e_1599 = {_e_1600, _e_1601};
    assign _e_1603 = 178;
    assign _e_1604 = 189;
    assign _e_1602 = {_e_1603, _e_1604};
    assign _e_1606 = 178;
    assign _e_1607 = 61;
    assign _e_1605 = {_e_1606, _e_1607};
    assign _e_1609 = 61;
    assign _e_1610 = 0;
    assign _e_1608 = {_e_1609, _e_1610};
    assign _e_1612 = 189;
    assign _e_1613 = 0;
    assign _e_1611 = {_e_1612, _e_1613};
    assign _e_1615 = 189;
    assign _e_1616 = 61;
    assign _e_1614 = {_e_1615, _e_1616};
    assign _e_1618 = 189;
    assign _e_1619 = 189;
    assign _e_1617 = {_e_1618, _e_1619};
    assign _e_1621 = 189;
    assign _e_1622 = 61;
    assign _e_1620 = {_e_1621, _e_1622};
    assign _e_1624 = 61;
    assign _e_1625 = 0;
    assign _e_1623 = {_e_1624, _e_1625};
    assign _e_1627 = 189;
    assign _e_1628 = 0;
    assign _e_1626 = {_e_1627, _e_1628};
    assign _e_1630 = 179;
    assign _e_1631 = 61;
    assign _e_1629 = {_e_1630, _e_1631};
    assign _e_1633 = 179;
    assign _e_1634 = 189;
    assign _e_1632 = {_e_1633, _e_1634};
    assign _e_1636 = 179;
    assign _e_1637 = 61;
    assign _e_1635 = {_e_1636, _e_1637};
    assign _e_1639 = 52;
    assign _e_1640 = 0;
    assign _e_1638 = {_e_1639, _e_1640};
    assign _e_1642 = 180;
    assign _e_1643 = 0;
    assign _e_1641 = {_e_1642, _e_1643};
    assign _e_1645 = 178;
    assign _e_1646 = 62;
    assign _e_1644 = {_e_1645, _e_1646};
    assign _e_1648 = 178;
    assign _e_1649 = 190;
    assign _e_1647 = {_e_1648, _e_1649};
    assign _e_1651 = 178;
    assign _e_1652 = 62;
    assign _e_1650 = {_e_1651, _e_1652};
    assign _e_1654 = 62;
    assign _e_1655 = 0;
    assign _e_1653 = {_e_1654, _e_1655};
    assign _e_1657 = 190;
    assign _e_1658 = 0;
    assign _e_1656 = {_e_1657, _e_1658};
    assign _e_1660 = 190;
    assign _e_1661 = 62;
    assign _e_1659 = {_e_1660, _e_1661};
    assign _e_1663 = 190;
    assign _e_1664 = 190;
    assign _e_1662 = {_e_1663, _e_1664};
    assign _e_1666 = 190;
    assign _e_1667 = 62;
    assign _e_1665 = {_e_1666, _e_1667};
    assign _e_1669 = 62;
    assign _e_1670 = 0;
    assign _e_1668 = {_e_1669, _e_1670};
    assign _e_1672 = 190;
    assign _e_1673 = 0;
    assign _e_1671 = {_e_1672, _e_1673};
    assign _e_1675 = 128;
    assign _e_1676 = 62;
    assign _e_1674 = {_e_1675, _e_1676};
    assign _e_1678 = 128;
    assign _e_1679 = 190;
    assign _e_1677 = {_e_1678, _e_1679};
    assign _e_1681 = 128;
    assign _e_1682 = 62;
    assign _e_1680 = {_e_1681, _e_1682};
    assign _e_1684 = 20;
    assign _e_1685 = 0;
    assign _e_1683 = {_e_1684, _e_1685};
    assign _e_1687 = 148;
    assign _e_1688 = 0;
    assign _e_1686 = {_e_1687, _e_1688};
    assign _e_1690 = 141;
    assign _e_1691 = 63;
    assign _e_1689 = {_e_1690, _e_1691};
    assign _e_1693 = 141;
    assign _e_1694 = 191;
    assign _e_1692 = {_e_1693, _e_1694};
    assign _e_1696 = 141;
    assign _e_1697 = 63;
    assign _e_1695 = {_e_1696, _e_1697};
    assign _e_1699 = 63;
    assign _e_1700 = 0;
    assign _e_1698 = {_e_1699, _e_1700};
    assign _e_1702 = 191;
    assign _e_1703 = 0;
    assign _e_1701 = {_e_1702, _e_1703};
    assign _e_1705 = 191;
    assign _e_1706 = 63;
    assign _e_1704 = {_e_1705, _e_1706};
    assign _e_1708 = 191;
    assign _e_1709 = 191;
    assign _e_1707 = {_e_1708, _e_1709};
    assign _e_1711 = 191;
    assign _e_1712 = 63;
    assign _e_1710 = {_e_1711, _e_1712};
    assign _e_1714 = 63;
    assign _e_1715 = 0;
    assign _e_1713 = {_e_1714, _e_1715};
    assign _e_1717 = 191;
    assign _e_1718 = 0;
    assign _e_1716 = {_e_1717, _e_1718};
    assign _e_1720 = 128;
    assign _e_1721 = 63;
    assign _e_1719 = {_e_1720, _e_1721};
    assign _e_1723 = 128;
    assign _e_1724 = 191;
    assign _e_1722 = {_e_1723, _e_1724};
    assign _e_1726 = 128;
    assign _e_1727 = 63;
    assign _e_1725 = {_e_1726, _e_1727};
    assign _e_1729 = 52;
    assign _e_1730 = 0;
    assign _e_1728 = {_e_1729, _e_1730};
    assign _e_1732 = 180;
    assign _e_1733 = 0;
    assign _e_1731 = {_e_1732, _e_1733};
    assign _e_1735 = 141;
    assign _e_1736 = 64;
    assign _e_1734 = {_e_1735, _e_1736};
    assign _e_1738 = 141;
    assign _e_1739 = 192;
    assign _e_1737 = {_e_1738, _e_1739};
    assign _e_1741 = 141;
    assign _e_1742 = 64;
    assign _e_1740 = {_e_1741, _e_1742};
    assign _e_1744 = 64;
    assign _e_1745 = 0;
    assign _e_1743 = {_e_1744, _e_1745};
    assign _e_1747 = 192;
    assign _e_1748 = 0;
    assign _e_1746 = {_e_1747, _e_1748};
    assign _e_1750 = 192;
    assign _e_1751 = 64;
    assign _e_1749 = {_e_1750, _e_1751};
    assign _e_1753 = 192;
    assign _e_1754 = 192;
    assign _e_1752 = {_e_1753, _e_1754};
    assign _e_1756 = 192;
    assign _e_1757 = 64;
    assign _e_1755 = {_e_1756, _e_1757};
    assign _e_1759 = 64;
    assign _e_1760 = 0;
    assign _e_1758 = {_e_1759, _e_1760};
    assign _e_1762 = 192;
    assign _e_1763 = 0;
    assign _e_1761 = {_e_1762, _e_1763};
    assign _e_1765 = 179;
    assign _e_1766 = 64;
    assign _e_1764 = {_e_1765, _e_1766};
    assign _e_1768 = 179;
    assign _e_1769 = 192;
    assign _e_1767 = {_e_1768, _e_1769};
    assign _e_1771 = 179;
    assign _e_1772 = 64;
    assign _e_1770 = {_e_1771, _e_1772};
    assign _e_1774 = 61;
    assign _e_1775 = 0;
    assign _e_1773 = {_e_1774, _e_1775};
    assign _e_1777 = 189;
    assign _e_1778 = 0;
    assign _e_1776 = {_e_1777, _e_1778};
    assign _e_1780 = 190;
    assign _e_1781 = 127;
    assign _e_1779 = {_e_1780, _e_1781};
    assign _e_1783 = 190;
    assign _e_1784 = 255;
    assign _e_1782 = {_e_1783, _e_1784};
    assign _e_1786 = 190;
    assign _e_1787 = 127;
    assign _e_1785 = {_e_1786, _e_1787};
    assign _e_1789 = 127;
    assign _e_1790 = 0;
    assign _e_1788 = {_e_1789, _e_1790};
    assign _e_1792 = 255;
    assign _e_1793 = 0;
    assign _e_1791 = {_e_1792, _e_1793};
    assign _e_1795 = 255;
    assign _e_1796 = 127;
    assign _e_1794 = {_e_1795, _e_1796};
    assign _e_1798 = 255;
    assign _e_1799 = 255;
    assign _e_1797 = {_e_1798, _e_1799};
    assign _e_1801 = 255;
    assign _e_1802 = 127;
    assign _e_1800 = {_e_1801, _e_1802};
    assign _e_1804 = 63;
    assign _e_1805 = 0;
    assign _e_1803 = {_e_1804, _e_1805};
    assign _e_1807 = 191;
    assign _e_1808 = 0;
    assign _e_1806 = {_e_1807, _e_1808};
    assign _e_1810 = 192;
    assign _e_1811 = 33;
    assign _e_1809 = {_e_1810, _e_1811};
    assign _e_1813 = 192;
    assign _e_1814 = 161;
    assign _e_1812 = {_e_1813, _e_1814};
    assign _e_1816 = 192;
    assign _e_1817 = 33;
    assign _e_1815 = {_e_1816, _e_1817};
    assign _e_1819 = 33;
    assign _e_1820 = 0;
    assign _e_1818 = {_e_1819, _e_1820};
    assign _e_1822 = 161;
    assign _e_1823 = 0;
    assign _e_1821 = {_e_1822, _e_1823};
    assign _e_1825 = 161;
    assign _e_1826 = 33;
    assign _e_1824 = {_e_1825, _e_1826};
    assign _e_1828 = 161;
    assign _e_1829 = 161;
    assign _e_1827 = {_e_1828, _e_1829};
    assign _e_1831 = 161;
    assign _e_1832 = 33;
    assign _e_1830 = {_e_1831, _e_1832};
    assign _e_1834 = 33;
    assign _e_1835 = 0;
    assign _e_1833 = {_e_1834, _e_1835};
    assign _e_1837 = 161;
    assign _e_1838 = 0;
    assign _e_1836 = {_e_1837, _e_1838};
    assign _e_1840 = 255;
    assign _e_1841 = 33;
    assign _e_1839 = {_e_1840, _e_1841};
    assign _e_1843 = 255;
    assign _e_1844 = 161;
    assign _e_1842 = {_e_1843, _e_1844};
    assign _e_1846 = 255;
    assign _e_1847 = 33;
    assign _e_1845 = {_e_1846, _e_1847};
    assign _e_1849 = 13;
    assign _e_1850 = 0;
    assign _e_1848 = {_e_1849, _e_1850};
    assign _e_1852 = 141;
    assign _e_1853 = 0;
    assign _e_1851 = {_e_1852, _e_1853};
    assign _e_1855 = 128;
    assign _e_1856 = 61;
    assign _e_1854 = {_e_1855, _e_1856};
    assign _e_1858 = 128;
    assign _e_1859 = 189;
    assign _e_1857 = {_e_1858, _e_1859};
    assign _e_1861 = 128;
    assign _e_1862 = 61;
    assign _e_1860 = {_e_1861, _e_1862};
    assign _e_1864 = 20;
    assign _e_1865 = 0;
    assign _e_1863 = {_e_1864, _e_1865};
    assign _e_1867 = 148;
    assign _e_1868 = 0;
    assign _e_1866 = {_e_1867, _e_1868};
    assign _e_1870 = 141;
    assign _e_1871 = 62;
    assign _e_1869 = {_e_1870, _e_1871};
    assign _e_1873 = 141;
    assign _e_1874 = 190;
    assign _e_1872 = {_e_1873, _e_1874};
    assign _e_1876 = 141;
    assign _e_1877 = 62;
    assign _e_1875 = {_e_1876, _e_1877};
    assign _e_1879 = 20;
    assign _e_1880 = 0;
    assign _e_1878 = {_e_1879, _e_1880};
    assign _e_1882 = 148;
    assign _e_1883 = 0;
    assign _e_1881 = {_e_1882, _e_1883};
    assign _e_1885 = 128;
    assign _e_1886 = 63;
    assign _e_1884 = {_e_1885, _e_1886};
    assign _e_1888 = 128;
    assign _e_1889 = 191;
    assign _e_1887 = {_e_1888, _e_1889};
    assign _e_1891 = 128;
    assign _e_1892 = 63;
    assign _e_1890 = {_e_1891, _e_1892};
    assign _e_1894 = 61;
    assign _e_1895 = 0;
    assign _e_1893 = {_e_1894, _e_1895};
    assign _e_1897 = 189;
    assign _e_1898 = 0;
    assign _e_1896 = {_e_1897, _e_1898};
    assign _e_1900 = 190;
    assign _e_1901 = 20;
    assign _e_1899 = {_e_1900, _e_1901};
    assign _e_1903 = 190;
    assign _e_1904 = 148;
    assign _e_1902 = {_e_1903, _e_1904};
    assign _e_1906 = 190;
    assign _e_1907 = 20;
    assign _e_1905 = {_e_1906, _e_1907};
    assign _e_1909 = 20;
    assign _e_1910 = 0;
    assign _e_1908 = {_e_1909, _e_1910};
    assign _e_1912 = 148;
    assign _e_1913 = 0;
    assign _e_1911 = {_e_1912, _e_1913};
    assign _e_1915 = 148;
    assign _e_1916 = 20;
    assign _e_1914 = {_e_1915, _e_1916};
    assign _e_1918 = 148;
    assign _e_1919 = 148;
    assign _e_1917 = {_e_1918, _e_1919};
    assign _e_1921 = 148;
    assign _e_1922 = 20;
    assign _e_1920 = {_e_1921, _e_1922};
    assign _e_1924 = 20;
    assign _e_1925 = 0;
    assign _e_1923 = {_e_1924, _e_1925};
    assign _e_1927 = 148;
    assign _e_1928 = 0;
    assign _e_1926 = {_e_1927, _e_1928};
    assign _e_1930 = 191;
    assign _e_1931 = 20;
    assign _e_1929 = {_e_1930, _e_1931};
    assign _e_1933 = 191;
    assign _e_1934 = 148;
    assign _e_1932 = {_e_1933, _e_1934};
    assign _e_1936 = 191;
    assign _e_1937 = 20;
    assign _e_1935 = {_e_1936, _e_1937};
    assign _e_1939 = 14;
    assign _e_1940 = 0;
    assign _e_1938 = {_e_1939, _e_1940};
    assign _e_1942 = 142;
    assign _e_1943 = 0;
    assign _e_1941 = {_e_1942, _e_1943};
    assign _e_1945 = 142;
    assign _e_1946 = 50;
    assign _e_1944 = {_e_1945, _e_1946};
    assign _e_1948 = 142;
    assign _e_1949 = 178;
    assign _e_1947 = {_e_1948, _e_1949};
    assign _e_1951 = 142;
    assign _e_1952 = 50;
    assign _e_1950 = {_e_1951, _e_1952};
    assign _e_1954 = 0;
    assign _e_1955 = 0;
    assign _e_1953 = {_e_1954, _e_1955};
    assign _e_1957 = 128;
    assign _e_1958 = 0;
    assign _e_1956 = {_e_1957, _e_1958};
    assign _e_1960 = 128;
    assign _e_1961 = 51;
    assign _e_1959 = {_e_1960, _e_1961};
    assign _e_1963 = 128;
    assign _e_1964 = 179;
    assign _e_1962 = {_e_1963, _e_1964};
    assign _e_1966 = 128;
    assign _e_1967 = 51;
    assign _e_1965 = {_e_1966, _e_1967};
    assign _e_1969 = 20;
    assign _e_1970 = 0;
    assign _e_1968 = {_e_1969, _e_1970};
    assign _e_1972 = 148;
    assign _e_1973 = 0;
    assign _e_1971 = {_e_1972, _e_1973};
    assign _e_1975 = 148;
    assign _e_1976 = 52;
    assign _e_1974 = {_e_1975, _e_1976};
    assign _e_1978 = 148;
    assign _e_1979 = 180;
    assign _e_1977 = {_e_1978, _e_1979};
    assign _e_1981 = 148;
    assign _e_1982 = 52;
    assign _e_1980 = {_e_1981, _e_1982};
    assign _e_1984 = 20;
    assign _e_1985 = 0;
    assign _e_1983 = {_e_1984, _e_1985};
    assign _e_1987 = 148;
    assign _e_1988 = 0;
    assign _e_1986 = {_e_1987, _e_1988};
    assign _e_1990 = 178;
    assign _e_1991 = 61;
    assign _e_1989 = {_e_1990, _e_1991};
    assign _e_1993 = 178;
    assign _e_1994 = 189;
    assign _e_1992 = {_e_1993, _e_1994};
    assign _e_1996 = 178;
    assign _e_1997 = 61;
    assign _e_1995 = {_e_1996, _e_1997};
    assign _e_1999 = 61;
    assign _e_2000 = 0;
    assign _e_1998 = {_e_1999, _e_2000};
    assign _e_2002 = 189;
    assign _e_2003 = 0;
    assign _e_2001 = {_e_2002, _e_2003};
    assign _e_2005 = 189;
    assign _e_2006 = 61;
    assign _e_2004 = {_e_2005, _e_2006};
    assign _e_2008 = 189;
    assign _e_2009 = 189;
    assign _e_2007 = {_e_2008, _e_2009};
    assign _e_2011 = 189;
    assign _e_2012 = 61;
    assign _e_2010 = {_e_2011, _e_2012};
    assign _e_2014 = 61;
    assign _e_2015 = 0;
    assign _e_2013 = {_e_2014, _e_2015};
    assign _e_2017 = 189;
    assign _e_2018 = 0;
    assign _e_2016 = {_e_2017, _e_2018};
    assign _e_2020 = 179;
    assign _e_2021 = 61;
    assign _e_2019 = {_e_2020, _e_2021};
    assign _e_2023 = 179;
    assign _e_2024 = 189;
    assign _e_2022 = {_e_2023, _e_2024};
    assign _e_2026 = 179;
    assign _e_2027 = 61;
    assign _e_2025 = {_e_2026, _e_2027};
    assign _e_2029 = 52;
    assign _e_2030 = 0;
    assign _e_2028 = {_e_2029, _e_2030};
    assign _e_2032 = 180;
    assign _e_2033 = 0;
    assign _e_2031 = {_e_2032, _e_2033};
    assign _e_2035 = 178;
    assign _e_2036 = 62;
    assign _e_2034 = {_e_2035, _e_2036};
    assign _e_2038 = 178;
    assign _e_2039 = 190;
    assign _e_2037 = {_e_2038, _e_2039};
    assign _e_2041 = 178;
    assign _e_2042 = 62;
    assign _e_2040 = {_e_2041, _e_2042};
    assign _e_2044 = 62;
    assign _e_2045 = 0;
    assign _e_2043 = {_e_2044, _e_2045};
    assign _e_2047 = 190;
    assign _e_2048 = 0;
    assign _e_2046 = {_e_2047, _e_2048};
    assign _e_2050 = 190;
    assign _e_2051 = 62;
    assign _e_2049 = {_e_2050, _e_2051};
    assign _e_2053 = 190;
    assign _e_2054 = 190;
    assign _e_2052 = {_e_2053, _e_2054};
    assign _e_2056 = 190;
    assign _e_2057 = 62;
    assign _e_2055 = {_e_2056, _e_2057};
    assign _e_2059 = 62;
    assign _e_2060 = 0;
    assign _e_2058 = {_e_2059, _e_2060};
    assign _e_2062 = 190;
    assign _e_2063 = 0;
    assign _e_2061 = {_e_2062, _e_2063};
    assign _e_2065 = 128;
    assign _e_2066 = 62;
    assign _e_2064 = {_e_2065, _e_2066};
    assign _e_2068 = 128;
    assign _e_2069 = 190;
    assign _e_2067 = {_e_2068, _e_2069};
    assign _e_2071 = 128;
    assign _e_2072 = 62;
    assign _e_2070 = {_e_2071, _e_2072};
    assign _e_2074 = 20;
    assign _e_2075 = 0;
    assign _e_2073 = {_e_2074, _e_2075};
    assign _e_2077 = 148;
    assign _e_2078 = 0;
    assign _e_2076 = {_e_2077, _e_2078};
    assign _e_2080 = 142;
    assign _e_2081 = 63;
    assign _e_2079 = {_e_2080, _e_2081};
    assign _e_2083 = 142;
    assign _e_2084 = 191;
    assign _e_2082 = {_e_2083, _e_2084};
    assign _e_2086 = 142;
    assign _e_2087 = 63;
    assign _e_2085 = {_e_2086, _e_2087};
    assign _e_2089 = 63;
    assign _e_2090 = 0;
    assign _e_2088 = {_e_2089, _e_2090};
    assign _e_2092 = 191;
    assign _e_2093 = 0;
    assign _e_2091 = {_e_2092, _e_2093};
    assign _e_2095 = 191;
    assign _e_2096 = 63;
    assign _e_2094 = {_e_2095, _e_2096};
    assign _e_2098 = 191;
    assign _e_2099 = 191;
    assign _e_2097 = {_e_2098, _e_2099};
    assign _e_2101 = 191;
    assign _e_2102 = 63;
    assign _e_2100 = {_e_2101, _e_2102};
    assign _e_2104 = 63;
    assign _e_2105 = 0;
    assign _e_2103 = {_e_2104, _e_2105};
    assign _e_2107 = 191;
    assign _e_2108 = 0;
    assign _e_2106 = {_e_2107, _e_2108};
    assign _e_2110 = 128;
    assign _e_2111 = 63;
    assign _e_2109 = {_e_2110, _e_2111};
    assign _e_2113 = 128;
    assign _e_2114 = 191;
    assign _e_2112 = {_e_2113, _e_2114};
    assign _e_2116 = 128;
    assign _e_2117 = 63;
    assign _e_2115 = {_e_2116, _e_2117};
    assign _e_2119 = 52;
    assign _e_2120 = 0;
    assign _e_2118 = {_e_2119, _e_2120};
    assign _e_2122 = 180;
    assign _e_2123 = 0;
    assign _e_2121 = {_e_2122, _e_2123};
    assign _e_2125 = 142;
    assign _e_2126 = 64;
    assign _e_2124 = {_e_2125, _e_2126};
    assign _e_2128 = 142;
    assign _e_2129 = 192;
    assign _e_2127 = {_e_2128, _e_2129};
    assign _e_2131 = 142;
    assign _e_2132 = 64;
    assign _e_2130 = {_e_2131, _e_2132};
    assign _e_2134 = 64;
    assign _e_2135 = 0;
    assign _e_2133 = {_e_2134, _e_2135};
    assign _e_2137 = 192;
    assign _e_2138 = 0;
    assign _e_2136 = {_e_2137, _e_2138};
    assign _e_2140 = 192;
    assign _e_2141 = 64;
    assign _e_2139 = {_e_2140, _e_2141};
    assign _e_2143 = 192;
    assign _e_2144 = 192;
    assign _e_2142 = {_e_2143, _e_2144};
    assign _e_2146 = 192;
    assign _e_2147 = 64;
    assign _e_2145 = {_e_2146, _e_2147};
    assign _e_2149 = 64;
    assign _e_2150 = 0;
    assign _e_2148 = {_e_2149, _e_2150};
    assign _e_2152 = 192;
    assign _e_2153 = 0;
    assign _e_2151 = {_e_2152, _e_2153};
    assign _e_2155 = 179;
    assign _e_2156 = 64;
    assign _e_2154 = {_e_2155, _e_2156};
    assign _e_2158 = 179;
    assign _e_2159 = 192;
    assign _e_2157 = {_e_2158, _e_2159};
    assign _e_2161 = 179;
    assign _e_2162 = 64;
    assign _e_2160 = {_e_2161, _e_2162};
    assign _e_2164 = 61;
    assign _e_2165 = 0;
    assign _e_2163 = {_e_2164, _e_2165};
    assign _e_2167 = 189;
    assign _e_2168 = 0;
    assign _e_2166 = {_e_2167, _e_2168};
    assign _e_2170 = 190;
    assign _e_2171 = 127;
    assign _e_2169 = {_e_2170, _e_2171};
    assign _e_2173 = 190;
    assign _e_2174 = 255;
    assign _e_2172 = {_e_2173, _e_2174};
    assign _e_2176 = 190;
    assign _e_2177 = 127;
    assign _e_2175 = {_e_2176, _e_2177};
    assign _e_2179 = 127;
    assign _e_2180 = 0;
    assign _e_2178 = {_e_2179, _e_2180};
    assign _e_2182 = 255;
    assign _e_2183 = 0;
    assign _e_2181 = {_e_2182, _e_2183};
    assign _e_2185 = 255;
    assign _e_2186 = 127;
    assign _e_2184 = {_e_2185, _e_2186};
    assign _e_2188 = 255;
    assign _e_2189 = 255;
    assign _e_2187 = {_e_2188, _e_2189};
    assign _e_2191 = 255;
    assign _e_2192 = 127;
    assign _e_2190 = {_e_2191, _e_2192};
    assign _e_2194 = 63;
    assign _e_2195 = 0;
    assign _e_2193 = {_e_2194, _e_2195};
    assign _e_2197 = 191;
    assign _e_2198 = 0;
    assign _e_2196 = {_e_2197, _e_2198};
    assign _e_2200 = 192;
    assign _e_2201 = 34;
    assign _e_2199 = {_e_2200, _e_2201};
    assign _e_2203 = 192;
    assign _e_2204 = 162;
    assign _e_2202 = {_e_2203, _e_2204};
    assign _e_2206 = 192;
    assign _e_2207 = 34;
    assign _e_2205 = {_e_2206, _e_2207};
    assign _e_2209 = 34;
    assign _e_2210 = 0;
    assign _e_2208 = {_e_2209, _e_2210};
    assign _e_2212 = 162;
    assign _e_2213 = 0;
    assign _e_2211 = {_e_2212, _e_2213};
    assign _e_2215 = 162;
    assign _e_2216 = 34;
    assign _e_2214 = {_e_2215, _e_2216};
    assign _e_2218 = 162;
    assign _e_2219 = 162;
    assign _e_2217 = {_e_2218, _e_2219};
    assign _e_2221 = 162;
    assign _e_2222 = 34;
    assign _e_2220 = {_e_2221, _e_2222};
    assign _e_2224 = 34;
    assign _e_2225 = 0;
    assign _e_2223 = {_e_2224, _e_2225};
    assign _e_2227 = 162;
    assign _e_2228 = 0;
    assign _e_2226 = {_e_2227, _e_2228};
    assign _e_2230 = 255;
    assign _e_2231 = 34;
    assign _e_2229 = {_e_2230, _e_2231};
    assign _e_2233 = 255;
    assign _e_2234 = 162;
    assign _e_2232 = {_e_2233, _e_2234};
    assign _e_2236 = 255;
    assign _e_2237 = 34;
    assign _e_2235 = {_e_2236, _e_2237};
    assign _e_2239 = 14;
    assign _e_2240 = 0;
    assign _e_2238 = {_e_2239, _e_2240};
    assign _e_2242 = 142;
    assign _e_2243 = 0;
    assign _e_2241 = {_e_2242, _e_2243};
    assign _e_2245 = 128;
    assign _e_2246 = 61;
    assign _e_2244 = {_e_2245, _e_2246};
    assign _e_2248 = 128;
    assign _e_2249 = 189;
    assign _e_2247 = {_e_2248, _e_2249};
    assign _e_2251 = 128;
    assign _e_2252 = 61;
    assign _e_2250 = {_e_2251, _e_2252};
    assign _e_2254 = 20;
    assign _e_2255 = 0;
    assign _e_2253 = {_e_2254, _e_2255};
    assign _e_2257 = 148;
    assign _e_2258 = 0;
    assign _e_2256 = {_e_2257, _e_2258};
    assign _e_2260 = 142;
    assign _e_2261 = 62;
    assign _e_2259 = {_e_2260, _e_2261};
    assign _e_2263 = 142;
    assign _e_2264 = 190;
    assign _e_2262 = {_e_2263, _e_2264};
    assign _e_2266 = 142;
    assign _e_2267 = 62;
    assign _e_2265 = {_e_2266, _e_2267};
    assign _e_2269 = 20;
    assign _e_2270 = 0;
    assign _e_2268 = {_e_2269, _e_2270};
    assign _e_2272 = 148;
    assign _e_2273 = 0;
    assign _e_2271 = {_e_2272, _e_2273};
    assign _e_2275 = 128;
    assign _e_2276 = 63;
    assign _e_2274 = {_e_2275, _e_2276};
    assign _e_2278 = 128;
    assign _e_2279 = 191;
    assign _e_2277 = {_e_2278, _e_2279};
    assign _e_2281 = 128;
    assign _e_2282 = 63;
    assign _e_2280 = {_e_2281, _e_2282};
    assign _e_2284 = 61;
    assign _e_2285 = 0;
    assign _e_2283 = {_e_2284, _e_2285};
    assign _e_2287 = 189;
    assign _e_2288 = 0;
    assign _e_2286 = {_e_2287, _e_2288};
    assign _e_2290 = 190;
    assign _e_2291 = 20;
    assign _e_2289 = {_e_2290, _e_2291};
    assign _e_2293 = 190;
    assign _e_2294 = 148;
    assign _e_2292 = {_e_2293, _e_2294};
    assign _e_2296 = 190;
    assign _e_2297 = 20;
    assign _e_2295 = {_e_2296, _e_2297};
    assign _e_2299 = 20;
    assign _e_2300 = 0;
    assign _e_2298 = {_e_2299, _e_2300};
    assign _e_2302 = 148;
    assign _e_2303 = 0;
    assign _e_2301 = {_e_2302, _e_2303};
    assign _e_2305 = 148;
    assign _e_2306 = 20;
    assign _e_2304 = {_e_2305, _e_2306};
    assign _e_2308 = 148;
    assign _e_2309 = 148;
    assign _e_2307 = {_e_2308, _e_2309};
    assign _e_2311 = 148;
    assign _e_2312 = 20;
    assign _e_2310 = {_e_2311, _e_2312};
    assign _e_2314 = 20;
    assign _e_2315 = 0;
    assign _e_2313 = {_e_2314, _e_2315};
    assign _e_2317 = 148;
    assign _e_2318 = 0;
    assign _e_2316 = {_e_2317, _e_2318};
    assign _e_2320 = 191;
    assign _e_2321 = 20;
    assign _e_2319 = {_e_2320, _e_2321};
    assign _e_2323 = 191;
    assign _e_2324 = 148;
    assign _e_2322 = {_e_2323, _e_2324};
    assign _e_2326 = 191;
    assign _e_2327 = 20;
    assign _e_2325 = {_e_2326, _e_2327};
    assign _e_2329 = 15;
    assign _e_2330 = 0;
    assign _e_2328 = {_e_2329, _e_2330};
    assign _e_2332 = 143;
    assign _e_2333 = 0;
    assign _e_2331 = {_e_2332, _e_2333};
    assign _e_2335 = 143;
    assign _e_2336 = 50;
    assign _e_2334 = {_e_2335, _e_2336};
    assign _e_2338 = 143;
    assign _e_2339 = 178;
    assign _e_2337 = {_e_2338, _e_2339};
    assign _e_2341 = 143;
    assign _e_2342 = 50;
    assign _e_2340 = {_e_2341, _e_2342};
    assign _e_2344 = 0;
    assign _e_2345 = 0;
    assign _e_2343 = {_e_2344, _e_2345};
    assign _e_2347 = 128;
    assign _e_2348 = 0;
    assign _e_2346 = {_e_2347, _e_2348};
    assign _e_2350 = 128;
    assign _e_2351 = 51;
    assign _e_2349 = {_e_2350, _e_2351};
    assign _e_2353 = 128;
    assign _e_2354 = 179;
    assign _e_2352 = {_e_2353, _e_2354};
    assign _e_2356 = 128;
    assign _e_2357 = 51;
    assign _e_2355 = {_e_2356, _e_2357};
    assign _e_2359 = 20;
    assign _e_2360 = 0;
    assign _e_2358 = {_e_2359, _e_2360};
    assign _e_2362 = 148;
    assign _e_2363 = 0;
    assign _e_2361 = {_e_2362, _e_2363};
    assign _e_2365 = 148;
    assign _e_2366 = 52;
    assign _e_2364 = {_e_2365, _e_2366};
    assign _e_2368 = 148;
    assign _e_2369 = 180;
    assign _e_2367 = {_e_2368, _e_2369};
    assign _e_2371 = 148;
    assign _e_2372 = 52;
    assign _e_2370 = {_e_2371, _e_2372};
    assign _e_2374 = 20;
    assign _e_2375 = 0;
    assign _e_2373 = {_e_2374, _e_2375};
    assign _e_2377 = 148;
    assign _e_2378 = 0;
    assign _e_2376 = {_e_2377, _e_2378};
    assign _e_2380 = 178;
    assign _e_2381 = 61;
    assign _e_2379 = {_e_2380, _e_2381};
    assign _e_2383 = 178;
    assign _e_2384 = 189;
    assign _e_2382 = {_e_2383, _e_2384};
    assign _e_2386 = 178;
    assign _e_2387 = 61;
    assign _e_2385 = {_e_2386, _e_2387};
    assign _e_2389 = 61;
    assign _e_2390 = 0;
    assign _e_2388 = {_e_2389, _e_2390};
    assign _e_2392 = 189;
    assign _e_2393 = 0;
    assign _e_2391 = {_e_2392, _e_2393};
    assign _e_2395 = 189;
    assign _e_2396 = 61;
    assign _e_2394 = {_e_2395, _e_2396};
    assign _e_2398 = 189;
    assign _e_2399 = 189;
    assign _e_2397 = {_e_2398, _e_2399};
    assign _e_2401 = 189;
    assign _e_2402 = 61;
    assign _e_2400 = {_e_2401, _e_2402};
    assign _e_2404 = 61;
    assign _e_2405 = 0;
    assign _e_2403 = {_e_2404, _e_2405};
    assign _e_2407 = 189;
    assign _e_2408 = 0;
    assign _e_2406 = {_e_2407, _e_2408};
    assign _e_2410 = 179;
    assign _e_2411 = 61;
    assign _e_2409 = {_e_2410, _e_2411};
    assign _e_2413 = 179;
    assign _e_2414 = 189;
    assign _e_2412 = {_e_2413, _e_2414};
    assign _e_2416 = 179;
    assign _e_2417 = 61;
    assign _e_2415 = {_e_2416, _e_2417};
    assign _e_2419 = 52;
    assign _e_2420 = 0;
    assign _e_2418 = {_e_2419, _e_2420};
    assign _e_2422 = 180;
    assign _e_2423 = 0;
    assign _e_2421 = {_e_2422, _e_2423};
    assign _e_2425 = 178;
    assign _e_2426 = 62;
    assign _e_2424 = {_e_2425, _e_2426};
    assign _e_2428 = 178;
    assign _e_2429 = 190;
    assign _e_2427 = {_e_2428, _e_2429};
    assign _e_2431 = 178;
    assign _e_2432 = 62;
    assign _e_2430 = {_e_2431, _e_2432};
    assign _e_2434 = 62;
    assign _e_2435 = 0;
    assign _e_2433 = {_e_2434, _e_2435};
    assign _e_2437 = 190;
    assign _e_2438 = 0;
    assign _e_2436 = {_e_2437, _e_2438};
    assign _e_2440 = 190;
    assign _e_2441 = 62;
    assign _e_2439 = {_e_2440, _e_2441};
    assign _e_2443 = 190;
    assign _e_2444 = 190;
    assign _e_2442 = {_e_2443, _e_2444};
    assign _e_2446 = 190;
    assign _e_2447 = 62;
    assign _e_2445 = {_e_2446, _e_2447};
    assign _e_2449 = 62;
    assign _e_2450 = 0;
    assign _e_2448 = {_e_2449, _e_2450};
    assign _e_2452 = 190;
    assign _e_2453 = 0;
    assign _e_2451 = {_e_2452, _e_2453};
    assign _e_2455 = 128;
    assign _e_2456 = 62;
    assign _e_2454 = {_e_2455, _e_2456};
    assign _e_2458 = 128;
    assign _e_2459 = 190;
    assign _e_2457 = {_e_2458, _e_2459};
    assign _e_2461 = 128;
    assign _e_2462 = 62;
    assign _e_2460 = {_e_2461, _e_2462};
    assign _e_2464 = 20;
    assign _e_2465 = 0;
    assign _e_2463 = {_e_2464, _e_2465};
    assign _e_2467 = 148;
    assign _e_2468 = 0;
    assign _e_2466 = {_e_2467, _e_2468};
    assign _e_2470 = 143;
    assign _e_2471 = 63;
    assign _e_2469 = {_e_2470, _e_2471};
    assign _e_2473 = 143;
    assign _e_2474 = 191;
    assign _e_2472 = {_e_2473, _e_2474};
    assign _e_2476 = 143;
    assign _e_2477 = 63;
    assign _e_2475 = {_e_2476, _e_2477};
    assign _e_2479 = 63;
    assign _e_2480 = 0;
    assign _e_2478 = {_e_2479, _e_2480};
    assign _e_2482 = 191;
    assign _e_2483 = 0;
    assign _e_2481 = {_e_2482, _e_2483};
    assign _e_2485 = 191;
    assign _e_2486 = 63;
    assign _e_2484 = {_e_2485, _e_2486};
    assign _e_2488 = 191;
    assign _e_2489 = 191;
    assign _e_2487 = {_e_2488, _e_2489};
    assign _e_2491 = 191;
    assign _e_2492 = 63;
    assign _e_2490 = {_e_2491, _e_2492};
    assign _e_2494 = 63;
    assign _e_2495 = 0;
    assign _e_2493 = {_e_2494, _e_2495};
    assign _e_2497 = 191;
    assign _e_2498 = 0;
    assign _e_2496 = {_e_2497, _e_2498};
    assign _e_2500 = 128;
    assign _e_2501 = 63;
    assign _e_2499 = {_e_2500, _e_2501};
    assign _e_2503 = 128;
    assign _e_2504 = 191;
    assign _e_2502 = {_e_2503, _e_2504};
    assign _e_2506 = 128;
    assign _e_2507 = 63;
    assign _e_2505 = {_e_2506, _e_2507};
    assign _e_2509 = 52;
    assign _e_2510 = 0;
    assign _e_2508 = {_e_2509, _e_2510};
    assign _e_2512 = 180;
    assign _e_2513 = 0;
    assign _e_2511 = {_e_2512, _e_2513};
    assign _e_2515 = 143;
    assign _e_2516 = 64;
    assign _e_2514 = {_e_2515, _e_2516};
    assign _e_2518 = 143;
    assign _e_2519 = 192;
    assign _e_2517 = {_e_2518, _e_2519};
    assign _e_2521 = 143;
    assign _e_2522 = 64;
    assign _e_2520 = {_e_2521, _e_2522};
    assign _e_2524 = 64;
    assign _e_2525 = 0;
    assign _e_2523 = {_e_2524, _e_2525};
    assign _e_2527 = 192;
    assign _e_2528 = 0;
    assign _e_2526 = {_e_2527, _e_2528};
    assign _e_2530 = 192;
    assign _e_2531 = 64;
    assign _e_2529 = {_e_2530, _e_2531};
    assign _e_2533 = 192;
    assign _e_2534 = 192;
    assign _e_2532 = {_e_2533, _e_2534};
    assign _e_2536 = 192;
    assign _e_2537 = 64;
    assign _e_2535 = {_e_2536, _e_2537};
    assign _e_2539 = 64;
    assign _e_2540 = 0;
    assign _e_2538 = {_e_2539, _e_2540};
    assign _e_2542 = 192;
    assign _e_2543 = 0;
    assign _e_2541 = {_e_2542, _e_2543};
    assign _e_2545 = 179;
    assign _e_2546 = 64;
    assign _e_2544 = {_e_2545, _e_2546};
    assign _e_2548 = 179;
    assign _e_2549 = 192;
    assign _e_2547 = {_e_2548, _e_2549};
    assign _e_2551 = 179;
    assign _e_2552 = 64;
    assign _e_2550 = {_e_2551, _e_2552};
    assign _e_2554 = 61;
    assign _e_2555 = 0;
    assign _e_2553 = {_e_2554, _e_2555};
    assign _e_2557 = 189;
    assign _e_2558 = 0;
    assign _e_2556 = {_e_2557, _e_2558};
    assign _e_2560 = 190;
    assign _e_2561 = 127;
    assign _e_2559 = {_e_2560, _e_2561};
    assign _e_2563 = 190;
    assign _e_2564 = 255;
    assign _e_2562 = {_e_2563, _e_2564};
    assign _e_2566 = 190;
    assign _e_2567 = 127;
    assign _e_2565 = {_e_2566, _e_2567};
    assign _e_2569 = 127;
    assign _e_2570 = 0;
    assign _e_2568 = {_e_2569, _e_2570};
    assign _e_2572 = 255;
    assign _e_2573 = 0;
    assign _e_2571 = {_e_2572, _e_2573};
    assign _e_2575 = 255;
    assign _e_2576 = 127;
    assign _e_2574 = {_e_2575, _e_2576};
    assign _e_2578 = 255;
    assign _e_2579 = 255;
    assign _e_2577 = {_e_2578, _e_2579};
    assign _e_2581 = 255;
    assign _e_2582 = 127;
    assign _e_2580 = {_e_2581, _e_2582};
    assign _e_2584 = 63;
    assign _e_2585 = 0;
    assign _e_2583 = {_e_2584, _e_2585};
    assign _e_2587 = 191;
    assign _e_2588 = 0;
    assign _e_2586 = {_e_2587, _e_2588};
    assign _e_2590 = 192;
    assign _e_2591 = 35;
    assign _e_2589 = {_e_2590, _e_2591};
    assign _e_2593 = 192;
    assign _e_2594 = 163;
    assign _e_2592 = {_e_2593, _e_2594};
    assign _e_2596 = 192;
    assign _e_2597 = 35;
    assign _e_2595 = {_e_2596, _e_2597};
    assign _e_2599 = 35;
    assign _e_2600 = 0;
    assign _e_2598 = {_e_2599, _e_2600};
    assign _e_2602 = 163;
    assign _e_2603 = 0;
    assign _e_2601 = {_e_2602, _e_2603};
    assign _e_2605 = 163;
    assign _e_2606 = 35;
    assign _e_2604 = {_e_2605, _e_2606};
    assign _e_2608 = 163;
    assign _e_2609 = 163;
    assign _e_2607 = {_e_2608, _e_2609};
    assign _e_2611 = 163;
    assign _e_2612 = 35;
    assign _e_2610 = {_e_2611, _e_2612};
    assign _e_2614 = 35;
    assign _e_2615 = 0;
    assign _e_2613 = {_e_2614, _e_2615};
    assign _e_2617 = 163;
    assign _e_2618 = 0;
    assign _e_2616 = {_e_2617, _e_2618};
    assign _e_2620 = 255;
    assign _e_2621 = 35;
    assign _e_2619 = {_e_2620, _e_2621};
    assign _e_2623 = 255;
    assign _e_2624 = 163;
    assign _e_2622 = {_e_2623, _e_2624};
    assign _e_2626 = 255;
    assign _e_2627 = 35;
    assign _e_2625 = {_e_2626, _e_2627};
    assign _e_2629 = 15;
    assign _e_2630 = 0;
    assign _e_2628 = {_e_2629, _e_2630};
    assign _e_2632 = 143;
    assign _e_2633 = 0;
    assign _e_2631 = {_e_2632, _e_2633};
    assign _e_2635 = 128;
    assign _e_2636 = 61;
    assign _e_2634 = {_e_2635, _e_2636};
    assign _e_2638 = 128;
    assign _e_2639 = 189;
    assign _e_2637 = {_e_2638, _e_2639};
    assign _e_2641 = 128;
    assign _e_2642 = 61;
    assign _e_2640 = {_e_2641, _e_2642};
    assign _e_2644 = 20;
    assign _e_2645 = 0;
    assign _e_2643 = {_e_2644, _e_2645};
    assign _e_2647 = 148;
    assign _e_2648 = 0;
    assign _e_2646 = {_e_2647, _e_2648};
    assign _e_2650 = 143;
    assign _e_2651 = 62;
    assign _e_2649 = {_e_2650, _e_2651};
    assign _e_2653 = 143;
    assign _e_2654 = 190;
    assign _e_2652 = {_e_2653, _e_2654};
    assign _e_2656 = 143;
    assign _e_2657 = 62;
    assign _e_2655 = {_e_2656, _e_2657};
    assign _e_2659 = 20;
    assign _e_2660 = 0;
    assign _e_2658 = {_e_2659, _e_2660};
    assign _e_2662 = 148;
    assign _e_2663 = 0;
    assign _e_2661 = {_e_2662, _e_2663};
    assign _e_2665 = 128;
    assign _e_2666 = 63;
    assign _e_2664 = {_e_2665, _e_2666};
    assign _e_2668 = 128;
    assign _e_2669 = 191;
    assign _e_2667 = {_e_2668, _e_2669};
    assign _e_2671 = 128;
    assign _e_2672 = 63;
    assign _e_2670 = {_e_2671, _e_2672};
    assign _e_2674 = 61;
    assign _e_2675 = 0;
    assign _e_2673 = {_e_2674, _e_2675};
    assign _e_2677 = 189;
    assign _e_2678 = 0;
    assign _e_2676 = {_e_2677, _e_2678};
    assign _e_2680 = 190;
    assign _e_2681 = 20;
    assign _e_2679 = {_e_2680, _e_2681};
    assign _e_2683 = 190;
    assign _e_2684 = 148;
    assign _e_2682 = {_e_2683, _e_2684};
    assign _e_2686 = 190;
    assign _e_2687 = 20;
    assign _e_2685 = {_e_2686, _e_2687};
    assign _e_2689 = 20;
    assign _e_2690 = 0;
    assign _e_2688 = {_e_2689, _e_2690};
    assign _e_2692 = 148;
    assign _e_2693 = 0;
    assign _e_2691 = {_e_2692, _e_2693};
    assign _e_2695 = 148;
    assign _e_2696 = 20;
    assign _e_2694 = {_e_2695, _e_2696};
    assign _e_2698 = 148;
    assign _e_2699 = 148;
    assign _e_2697 = {_e_2698, _e_2699};
    assign _e_2701 = 148;
    assign _e_2702 = 20;
    assign _e_2700 = {_e_2701, _e_2702};
    assign _e_2704 = 20;
    assign _e_2705 = 0;
    assign _e_2703 = {_e_2704, _e_2705};
    assign _e_2707 = 148;
    assign _e_2708 = 0;
    assign _e_2706 = {_e_2707, _e_2708};
    assign _e_2710 = 191;
    assign _e_2711 = 20;
    assign _e_2709 = {_e_2710, _e_2711};
    assign _e_2713 = 191;
    assign _e_2714 = 148;
    assign _e_2712 = {_e_2713, _e_2714};
    assign _e_2716 = 191;
    assign _e_2717 = 20;
    assign _e_2715 = {_e_2716, _e_2717};
    assign _e_2719 = 16;
    assign _e_2720 = 0;
    assign _e_2718 = {_e_2719, _e_2720};
    assign _e_2722 = 144;
    assign _e_2723 = 0;
    assign _e_2721 = {_e_2722, _e_2723};
    assign _e_2725 = 144;
    assign _e_2726 = 50;
    assign _e_2724 = {_e_2725, _e_2726};
    assign _e_2728 = 144;
    assign _e_2729 = 178;
    assign _e_2727 = {_e_2728, _e_2729};
    assign _e_2731 = 144;
    assign _e_2732 = 50;
    assign _e_2730 = {_e_2731, _e_2732};
    assign _e_2734 = 0;
    assign _e_2735 = 0;
    assign _e_2733 = {_e_2734, _e_2735};
    assign _e_2737 = 128;
    assign _e_2738 = 0;
    assign _e_2736 = {_e_2737, _e_2738};
    assign _e_2740 = 128;
    assign _e_2741 = 51;
    assign _e_2739 = {_e_2740, _e_2741};
    assign _e_2743 = 128;
    assign _e_2744 = 179;
    assign _e_2742 = {_e_2743, _e_2744};
    assign _e_2746 = 128;
    assign _e_2747 = 51;
    assign _e_2745 = {_e_2746, _e_2747};
    assign _e_2749 = 20;
    assign _e_2750 = 0;
    assign _e_2748 = {_e_2749, _e_2750};
    assign _e_2752 = 148;
    assign _e_2753 = 0;
    assign _e_2751 = {_e_2752, _e_2753};
    assign _e_2755 = 148;
    assign _e_2756 = 52;
    assign _e_2754 = {_e_2755, _e_2756};
    assign _e_2758 = 148;
    assign _e_2759 = 180;
    assign _e_2757 = {_e_2758, _e_2759};
    assign _e_2761 = 148;
    assign _e_2762 = 52;
    assign _e_2760 = {_e_2761, _e_2762};
    assign _e_2764 = 20;
    assign _e_2765 = 0;
    assign _e_2763 = {_e_2764, _e_2765};
    assign _e_2767 = 148;
    assign _e_2768 = 0;
    assign _e_2766 = {_e_2767, _e_2768};
    assign _e_2770 = 178;
    assign _e_2771 = 61;
    assign _e_2769 = {_e_2770, _e_2771};
    assign _e_2773 = 178;
    assign _e_2774 = 189;
    assign _e_2772 = {_e_2773, _e_2774};
    assign _e_2776 = 178;
    assign _e_2777 = 61;
    assign _e_2775 = {_e_2776, _e_2777};
    assign _e_2779 = 61;
    assign _e_2780 = 0;
    assign _e_2778 = {_e_2779, _e_2780};
    assign _e_2782 = 189;
    assign _e_2783 = 0;
    assign _e_2781 = {_e_2782, _e_2783};
    assign _e_2785 = 189;
    assign _e_2786 = 61;
    assign _e_2784 = {_e_2785, _e_2786};
    assign _e_2788 = 189;
    assign _e_2789 = 189;
    assign _e_2787 = {_e_2788, _e_2789};
    assign _e_2791 = 189;
    assign _e_2792 = 61;
    assign _e_2790 = {_e_2791, _e_2792};
    assign _e_2794 = 61;
    assign _e_2795 = 0;
    assign _e_2793 = {_e_2794, _e_2795};
    assign _e_2797 = 189;
    assign _e_2798 = 0;
    assign _e_2796 = {_e_2797, _e_2798};
    assign _e_2800 = 179;
    assign _e_2801 = 61;
    assign _e_2799 = {_e_2800, _e_2801};
    assign _e_2803 = 179;
    assign _e_2804 = 189;
    assign _e_2802 = {_e_2803, _e_2804};
    assign _e_2806 = 179;
    assign _e_2807 = 61;
    assign _e_2805 = {_e_2806, _e_2807};
    assign _e_2809 = 52;
    assign _e_2810 = 0;
    assign _e_2808 = {_e_2809, _e_2810};
    assign _e_2812 = 180;
    assign _e_2813 = 0;
    assign _e_2811 = {_e_2812, _e_2813};
    assign _e_2815 = 178;
    assign _e_2816 = 62;
    assign _e_2814 = {_e_2815, _e_2816};
    assign _e_2818 = 178;
    assign _e_2819 = 190;
    assign _e_2817 = {_e_2818, _e_2819};
    assign _e_2821 = 178;
    assign _e_2822 = 62;
    assign _e_2820 = {_e_2821, _e_2822};
    assign _e_2824 = 62;
    assign _e_2825 = 0;
    assign _e_2823 = {_e_2824, _e_2825};
    assign _e_2827 = 190;
    assign _e_2828 = 0;
    assign _e_2826 = {_e_2827, _e_2828};
    assign _e_2830 = 190;
    assign _e_2831 = 62;
    assign _e_2829 = {_e_2830, _e_2831};
    assign _e_2833 = 190;
    assign _e_2834 = 190;
    assign _e_2832 = {_e_2833, _e_2834};
    assign _e_2836 = 190;
    assign _e_2837 = 62;
    assign _e_2835 = {_e_2836, _e_2837};
    assign _e_2839 = 62;
    assign _e_2840 = 0;
    assign _e_2838 = {_e_2839, _e_2840};
    assign _e_2842 = 190;
    assign _e_2843 = 0;
    assign _e_2841 = {_e_2842, _e_2843};
    assign _e_2845 = 128;
    assign _e_2846 = 62;
    assign _e_2844 = {_e_2845, _e_2846};
    assign _e_2848 = 128;
    assign _e_2849 = 190;
    assign _e_2847 = {_e_2848, _e_2849};
    assign _e_2851 = 128;
    assign _e_2852 = 62;
    assign _e_2850 = {_e_2851, _e_2852};
    assign _e_2854 = 20;
    assign _e_2855 = 0;
    assign _e_2853 = {_e_2854, _e_2855};
    assign _e_2857 = 148;
    assign _e_2858 = 0;
    assign _e_2856 = {_e_2857, _e_2858};
    assign _e_2860 = 144;
    assign _e_2861 = 63;
    assign _e_2859 = {_e_2860, _e_2861};
    assign _e_2863 = 144;
    assign _e_2864 = 191;
    assign _e_2862 = {_e_2863, _e_2864};
    assign _e_2866 = 144;
    assign _e_2867 = 63;
    assign _e_2865 = {_e_2866, _e_2867};
    assign _e_2869 = 63;
    assign _e_2870 = 0;
    assign _e_2868 = {_e_2869, _e_2870};
    assign _e_2872 = 191;
    assign _e_2873 = 0;
    assign _e_2871 = {_e_2872, _e_2873};
    assign _e_2875 = 191;
    assign _e_2876 = 63;
    assign _e_2874 = {_e_2875, _e_2876};
    assign _e_2878 = 191;
    assign _e_2879 = 191;
    assign _e_2877 = {_e_2878, _e_2879};
    assign _e_2881 = 191;
    assign _e_2882 = 63;
    assign _e_2880 = {_e_2881, _e_2882};
    assign _e_2884 = 63;
    assign _e_2885 = 0;
    assign _e_2883 = {_e_2884, _e_2885};
    assign _e_2887 = 191;
    assign _e_2888 = 0;
    assign _e_2886 = {_e_2887, _e_2888};
    assign _e_2890 = 128;
    assign _e_2891 = 63;
    assign _e_2889 = {_e_2890, _e_2891};
    assign _e_2893 = 128;
    assign _e_2894 = 191;
    assign _e_2892 = {_e_2893, _e_2894};
    assign _e_2896 = 128;
    assign _e_2897 = 63;
    assign _e_2895 = {_e_2896, _e_2897};
    assign _e_2899 = 52;
    assign _e_2900 = 0;
    assign _e_2898 = {_e_2899, _e_2900};
    assign _e_2902 = 180;
    assign _e_2903 = 0;
    assign _e_2901 = {_e_2902, _e_2903};
    assign _e_2905 = 144;
    assign _e_2906 = 64;
    assign _e_2904 = {_e_2905, _e_2906};
    assign _e_2908 = 144;
    assign _e_2909 = 192;
    assign _e_2907 = {_e_2908, _e_2909};
    assign _e_2911 = 144;
    assign _e_2912 = 64;
    assign _e_2910 = {_e_2911, _e_2912};
    assign _e_2914 = 64;
    assign _e_2915 = 0;
    assign _e_2913 = {_e_2914, _e_2915};
    assign _e_2917 = 192;
    assign _e_2918 = 0;
    assign _e_2916 = {_e_2917, _e_2918};
    assign _e_2920 = 192;
    assign _e_2921 = 64;
    assign _e_2919 = {_e_2920, _e_2921};
    assign _e_2923 = 192;
    assign _e_2924 = 192;
    assign _e_2922 = {_e_2923, _e_2924};
    assign _e_2926 = 192;
    assign _e_2927 = 64;
    assign _e_2925 = {_e_2926, _e_2927};
    assign _e_2929 = 64;
    assign _e_2930 = 0;
    assign _e_2928 = {_e_2929, _e_2930};
    assign _e_2932 = 192;
    assign _e_2933 = 0;
    assign _e_2931 = {_e_2932, _e_2933};
    assign _e_2935 = 179;
    assign _e_2936 = 64;
    assign _e_2934 = {_e_2935, _e_2936};
    assign _e_2938 = 179;
    assign _e_2939 = 192;
    assign _e_2937 = {_e_2938, _e_2939};
    assign _e_2941 = 179;
    assign _e_2942 = 64;
    assign _e_2940 = {_e_2941, _e_2942};
    assign _e_2944 = 61;
    assign _e_2945 = 0;
    assign _e_2943 = {_e_2944, _e_2945};
    assign _e_2947 = 189;
    assign _e_2948 = 0;
    assign _e_2946 = {_e_2947, _e_2948};
    assign _e_2950 = 190;
    assign _e_2951 = 127;
    assign _e_2949 = {_e_2950, _e_2951};
    assign _e_2953 = 190;
    assign _e_2954 = 255;
    assign _e_2952 = {_e_2953, _e_2954};
    assign _e_2956 = 190;
    assign _e_2957 = 127;
    assign _e_2955 = {_e_2956, _e_2957};
    assign _e_2959 = 127;
    assign _e_2960 = 0;
    assign _e_2958 = {_e_2959, _e_2960};
    assign _e_2962 = 255;
    assign _e_2963 = 0;
    assign _e_2961 = {_e_2962, _e_2963};
    assign _e_2965 = 255;
    assign _e_2966 = 127;
    assign _e_2964 = {_e_2965, _e_2966};
    assign _e_2968 = 255;
    assign _e_2969 = 255;
    assign _e_2967 = {_e_2968, _e_2969};
    assign _e_2971 = 255;
    assign _e_2972 = 127;
    assign _e_2970 = {_e_2971, _e_2972};
    assign _e_2974 = 63;
    assign _e_2975 = 0;
    assign _e_2973 = {_e_2974, _e_2975};
    assign _e_2977 = 191;
    assign _e_2978 = 0;
    assign _e_2976 = {_e_2977, _e_2978};
    assign _e_2980 = 192;
    assign _e_2981 = 36;
    assign _e_2979 = {_e_2980, _e_2981};
    assign _e_2983 = 192;
    assign _e_2984 = 164;
    assign _e_2982 = {_e_2983, _e_2984};
    assign _e_2986 = 192;
    assign _e_2987 = 36;
    assign _e_2985 = {_e_2986, _e_2987};
    assign _e_2989 = 36;
    assign _e_2990 = 0;
    assign _e_2988 = {_e_2989, _e_2990};
    assign _e_2992 = 164;
    assign _e_2993 = 0;
    assign _e_2991 = {_e_2992, _e_2993};
    assign _e_2995 = 164;
    assign _e_2996 = 36;
    assign _e_2994 = {_e_2995, _e_2996};
    assign _e_2998 = 164;
    assign _e_2999 = 164;
    assign _e_2997 = {_e_2998, _e_2999};
    assign _e_3001 = 164;
    assign _e_3002 = 36;
    assign _e_3000 = {_e_3001, _e_3002};
    assign _e_3004 = 36;
    assign _e_3005 = 0;
    assign _e_3003 = {_e_3004, _e_3005};
    assign _e_3007 = 164;
    assign _e_3008 = 0;
    assign _e_3006 = {_e_3007, _e_3008};
    assign _e_3010 = 255;
    assign _e_3011 = 36;
    assign _e_3009 = {_e_3010, _e_3011};
    assign _e_3013 = 255;
    assign _e_3014 = 164;
    assign _e_3012 = {_e_3013, _e_3014};
    assign _e_3016 = 255;
    assign _e_3017 = 36;
    assign _e_3015 = {_e_3016, _e_3017};
    assign _e_3019 = 16;
    assign _e_3020 = 0;
    assign _e_3018 = {_e_3019, _e_3020};
    assign _e_3022 = 144;
    assign _e_3023 = 0;
    assign _e_3021 = {_e_3022, _e_3023};
    assign _e_3025 = 128;
    assign _e_3026 = 61;
    assign _e_3024 = {_e_3025, _e_3026};
    assign _e_3028 = 128;
    assign _e_3029 = 189;
    assign _e_3027 = {_e_3028, _e_3029};
    assign _e_3031 = 128;
    assign _e_3032 = 61;
    assign _e_3030 = {_e_3031, _e_3032};
    assign _e_3034 = 20;
    assign _e_3035 = 0;
    assign _e_3033 = {_e_3034, _e_3035};
    assign _e_3037 = 148;
    assign _e_3038 = 0;
    assign _e_3036 = {_e_3037, _e_3038};
    assign _e_3040 = 144;
    assign _e_3041 = 62;
    assign _e_3039 = {_e_3040, _e_3041};
    assign _e_3043 = 144;
    assign _e_3044 = 190;
    assign _e_3042 = {_e_3043, _e_3044};
    assign _e_3046 = 144;
    assign _e_3047 = 62;
    assign _e_3045 = {_e_3046, _e_3047};
    assign _e_3049 = 20;
    assign _e_3050 = 0;
    assign _e_3048 = {_e_3049, _e_3050};
    assign _e_3052 = 148;
    assign _e_3053 = 0;
    assign _e_3051 = {_e_3052, _e_3053};
    assign _e_3055 = 128;
    assign _e_3056 = 63;
    assign _e_3054 = {_e_3055, _e_3056};
    assign _e_3058 = 128;
    assign _e_3059 = 191;
    assign _e_3057 = {_e_3058, _e_3059};
    assign _e_3061 = 128;
    assign _e_3062 = 63;
    assign _e_3060 = {_e_3061, _e_3062};
    assign _e_3064 = 61;
    assign _e_3065 = 0;
    assign _e_3063 = {_e_3064, _e_3065};
    assign _e_3067 = 189;
    assign _e_3068 = 0;
    assign _e_3066 = {_e_3067, _e_3068};
    assign _e_3070 = 190;
    assign _e_3071 = 20;
    assign _e_3069 = {_e_3070, _e_3071};
    assign _e_3073 = 190;
    assign _e_3074 = 148;
    assign _e_3072 = {_e_3073, _e_3074};
    assign _e_3076 = 190;
    assign _e_3077 = 20;
    assign _e_3075 = {_e_3076, _e_3077};
    assign _e_3079 = 20;
    assign _e_3080 = 0;
    assign _e_3078 = {_e_3079, _e_3080};
    assign _e_3082 = 148;
    assign _e_3083 = 0;
    assign _e_3081 = {_e_3082, _e_3083};
    assign _e_3085 = 148;
    assign _e_3086 = 20;
    assign _e_3084 = {_e_3085, _e_3086};
    assign _e_3088 = 148;
    assign _e_3089 = 148;
    assign _e_3087 = {_e_3088, _e_3089};
    assign _e_3091 = 148;
    assign _e_3092 = 20;
    assign _e_3090 = {_e_3091, _e_3092};
    assign _e_3094 = 20;
    assign _e_3095 = 0;
    assign _e_3093 = {_e_3094, _e_3095};
    assign _e_3097 = 148;
    assign _e_3098 = 0;
    assign _e_3096 = {_e_3097, _e_3098};
    assign _e_3100 = 191;
    assign _e_3101 = 20;
    assign _e_3099 = {_e_3100, _e_3101};
    assign _e_3103 = 191;
    assign _e_3104 = 148;
    assign _e_3102 = {_e_3103, _e_3104};
    assign _e_3106 = 191;
    assign _e_3107 = 20;
    assign _e_3105 = {_e_3106, _e_3107};
    assign _e_3109 = 17;
    assign _e_3110 = 0;
    assign _e_3108 = {_e_3109, _e_3110};
    assign _e_3112 = 145;
    assign _e_3113 = 0;
    assign _e_3111 = {_e_3112, _e_3113};
    assign _e_3115 = 145;
    assign _e_3116 = 50;
    assign _e_3114 = {_e_3115, _e_3116};
    assign _e_3118 = 145;
    assign _e_3119 = 178;
    assign _e_3117 = {_e_3118, _e_3119};
    assign _e_3121 = 145;
    assign _e_3122 = 50;
    assign _e_3120 = {_e_3121, _e_3122};
    assign _e_3124 = 0;
    assign _e_3125 = 0;
    assign _e_3123 = {_e_3124, _e_3125};
    assign _e_3127 = 128;
    assign _e_3128 = 0;
    assign _e_3126 = {_e_3127, _e_3128};
    assign _e_3130 = 128;
    assign _e_3131 = 51;
    assign _e_3129 = {_e_3130, _e_3131};
    assign _e_3133 = 128;
    assign _e_3134 = 179;
    assign _e_3132 = {_e_3133, _e_3134};
    assign _e_3136 = 128;
    assign _e_3137 = 51;
    assign _e_3135 = {_e_3136, _e_3137};
    assign _e_3139 = 20;
    assign _e_3140 = 0;
    assign _e_3138 = {_e_3139, _e_3140};
    assign _e_3142 = 148;
    assign _e_3143 = 0;
    assign _e_3141 = {_e_3142, _e_3143};
    assign _e_3145 = 148;
    assign _e_3146 = 52;
    assign _e_3144 = {_e_3145, _e_3146};
    assign _e_3148 = 148;
    assign _e_3149 = 180;
    assign _e_3147 = {_e_3148, _e_3149};
    assign _e_3151 = 148;
    assign _e_3152 = 52;
    assign _e_3150 = {_e_3151, _e_3152};
    assign _e_3154 = 20;
    assign _e_3155 = 0;
    assign _e_3153 = {_e_3154, _e_3155};
    assign _e_3157 = 148;
    assign _e_3158 = 0;
    assign _e_3156 = {_e_3157, _e_3158};
    assign _e_3160 = 178;
    assign _e_3161 = 61;
    assign _e_3159 = {_e_3160, _e_3161};
    assign _e_3163 = 178;
    assign _e_3164 = 189;
    assign _e_3162 = {_e_3163, _e_3164};
    assign _e_3166 = 178;
    assign _e_3167 = 61;
    assign _e_3165 = {_e_3166, _e_3167};
    assign _e_3169 = 61;
    assign _e_3170 = 0;
    assign _e_3168 = {_e_3169, _e_3170};
    assign _e_3172 = 189;
    assign _e_3173 = 0;
    assign _e_3171 = {_e_3172, _e_3173};
    assign _e_3175 = 189;
    assign _e_3176 = 61;
    assign _e_3174 = {_e_3175, _e_3176};
    assign _e_3178 = 189;
    assign _e_3179 = 189;
    assign _e_3177 = {_e_3178, _e_3179};
    assign _e_3181 = 189;
    assign _e_3182 = 61;
    assign _e_3180 = {_e_3181, _e_3182};
    assign _e_3184 = 61;
    assign _e_3185 = 0;
    assign _e_3183 = {_e_3184, _e_3185};
    assign _e_3187 = 189;
    assign _e_3188 = 0;
    assign _e_3186 = {_e_3187, _e_3188};
    assign _e_3190 = 179;
    assign _e_3191 = 61;
    assign _e_3189 = {_e_3190, _e_3191};
    assign _e_3193 = 179;
    assign _e_3194 = 189;
    assign _e_3192 = {_e_3193, _e_3194};
    assign _e_3196 = 179;
    assign _e_3197 = 61;
    assign _e_3195 = {_e_3196, _e_3197};
    assign _e_3199 = 52;
    assign _e_3200 = 0;
    assign _e_3198 = {_e_3199, _e_3200};
    assign _e_3202 = 180;
    assign _e_3203 = 0;
    assign _e_3201 = {_e_3202, _e_3203};
    assign _e_3205 = 178;
    assign _e_3206 = 62;
    assign _e_3204 = {_e_3205, _e_3206};
    assign _e_3208 = 178;
    assign _e_3209 = 190;
    assign _e_3207 = {_e_3208, _e_3209};
    assign _e_3211 = 178;
    assign _e_3212 = 62;
    assign _e_3210 = {_e_3211, _e_3212};
    assign _e_3214 = 62;
    assign _e_3215 = 0;
    assign _e_3213 = {_e_3214, _e_3215};
    assign _e_3217 = 190;
    assign _e_3218 = 0;
    assign _e_3216 = {_e_3217, _e_3218};
    assign _e_3220 = 190;
    assign _e_3221 = 62;
    assign _e_3219 = {_e_3220, _e_3221};
    assign _e_3223 = 190;
    assign _e_3224 = 190;
    assign _e_3222 = {_e_3223, _e_3224};
    assign _e_3226 = 190;
    assign _e_3227 = 62;
    assign _e_3225 = {_e_3226, _e_3227};
    assign _e_3229 = 62;
    assign _e_3230 = 0;
    assign _e_3228 = {_e_3229, _e_3230};
    assign _e_3232 = 190;
    assign _e_3233 = 0;
    assign _e_3231 = {_e_3232, _e_3233};
    assign _e_3235 = 128;
    assign _e_3236 = 62;
    assign _e_3234 = {_e_3235, _e_3236};
    assign _e_3238 = 128;
    assign _e_3239 = 190;
    assign _e_3237 = {_e_3238, _e_3239};
    assign _e_3241 = 128;
    assign _e_3242 = 62;
    assign _e_3240 = {_e_3241, _e_3242};
    assign _e_3244 = 20;
    assign _e_3245 = 0;
    assign _e_3243 = {_e_3244, _e_3245};
    assign _e_3247 = 148;
    assign _e_3248 = 0;
    assign _e_3246 = {_e_3247, _e_3248};
    assign _e_3250 = 145;
    assign _e_3251 = 63;
    assign _e_3249 = {_e_3250, _e_3251};
    assign _e_3253 = 145;
    assign _e_3254 = 191;
    assign _e_3252 = {_e_3253, _e_3254};
    assign _e_3256 = 145;
    assign _e_3257 = 63;
    assign _e_3255 = {_e_3256, _e_3257};
    assign _e_3259 = 63;
    assign _e_3260 = 0;
    assign _e_3258 = {_e_3259, _e_3260};
    assign _e_3262 = 191;
    assign _e_3263 = 0;
    assign _e_3261 = {_e_3262, _e_3263};
    assign _e_3265 = 191;
    assign _e_3266 = 63;
    assign _e_3264 = {_e_3265, _e_3266};
    assign _e_3268 = 191;
    assign _e_3269 = 191;
    assign _e_3267 = {_e_3268, _e_3269};
    assign _e_3271 = 191;
    assign _e_3272 = 63;
    assign _e_3270 = {_e_3271, _e_3272};
    assign _e_3274 = 63;
    assign _e_3275 = 0;
    assign _e_3273 = {_e_3274, _e_3275};
    assign _e_3277 = 191;
    assign _e_3278 = 0;
    assign _e_3276 = {_e_3277, _e_3278};
    assign _e_3280 = 128;
    assign _e_3281 = 63;
    assign _e_3279 = {_e_3280, _e_3281};
    assign _e_3283 = 128;
    assign _e_3284 = 191;
    assign _e_3282 = {_e_3283, _e_3284};
    assign _e_3286 = 128;
    assign _e_3287 = 63;
    assign _e_3285 = {_e_3286, _e_3287};
    assign _e_3289 = 52;
    assign _e_3290 = 0;
    assign _e_3288 = {_e_3289, _e_3290};
    assign _e_3292 = 180;
    assign _e_3293 = 0;
    assign _e_3291 = {_e_3292, _e_3293};
    assign _e_3295 = 145;
    assign _e_3296 = 64;
    assign _e_3294 = {_e_3295, _e_3296};
    assign _e_3298 = 145;
    assign _e_3299 = 192;
    assign _e_3297 = {_e_3298, _e_3299};
    assign _e_3301 = 145;
    assign _e_3302 = 64;
    assign _e_3300 = {_e_3301, _e_3302};
    assign _e_3304 = 64;
    assign _e_3305 = 0;
    assign _e_3303 = {_e_3304, _e_3305};
    assign _e_3307 = 192;
    assign _e_3308 = 0;
    assign _e_3306 = {_e_3307, _e_3308};
    assign _e_3310 = 192;
    assign _e_3311 = 64;
    assign _e_3309 = {_e_3310, _e_3311};
    assign _e_3313 = 192;
    assign _e_3314 = 192;
    assign _e_3312 = {_e_3313, _e_3314};
    assign _e_3316 = 192;
    assign _e_3317 = 64;
    assign _e_3315 = {_e_3316, _e_3317};
    assign _e_3319 = 64;
    assign _e_3320 = 0;
    assign _e_3318 = {_e_3319, _e_3320};
    assign _e_3322 = 192;
    assign _e_3323 = 0;
    assign _e_3321 = {_e_3322, _e_3323};
    assign _e_3325 = 179;
    assign _e_3326 = 64;
    assign _e_3324 = {_e_3325, _e_3326};
    assign _e_3328 = 179;
    assign _e_3329 = 192;
    assign _e_3327 = {_e_3328, _e_3329};
    assign _e_3331 = 179;
    assign _e_3332 = 64;
    assign _e_3330 = {_e_3331, _e_3332};
    assign _e_3334 = 61;
    assign _e_3335 = 0;
    assign _e_3333 = {_e_3334, _e_3335};
    assign _e_3337 = 189;
    assign _e_3338 = 0;
    assign _e_3336 = {_e_3337, _e_3338};
    assign _e_3340 = 190;
    assign _e_3341 = 127;
    assign _e_3339 = {_e_3340, _e_3341};
    assign _e_3343 = 190;
    assign _e_3344 = 255;
    assign _e_3342 = {_e_3343, _e_3344};
    assign _e_3346 = 190;
    assign _e_3347 = 127;
    assign _e_3345 = {_e_3346, _e_3347};
    assign _e_3349 = 127;
    assign _e_3350 = 0;
    assign _e_3348 = {_e_3349, _e_3350};
    assign _e_3352 = 255;
    assign _e_3353 = 0;
    assign _e_3351 = {_e_3352, _e_3353};
    assign _e_3355 = 255;
    assign _e_3356 = 127;
    assign _e_3354 = {_e_3355, _e_3356};
    assign _e_3358 = 255;
    assign _e_3359 = 255;
    assign _e_3357 = {_e_3358, _e_3359};
    assign _e_3361 = 255;
    assign _e_3362 = 127;
    assign _e_3360 = {_e_3361, _e_3362};
    assign _e_3364 = 63;
    assign _e_3365 = 0;
    assign _e_3363 = {_e_3364, _e_3365};
    assign _e_3367 = 191;
    assign _e_3368 = 0;
    assign _e_3366 = {_e_3367, _e_3368};
    assign _e_3370 = 192;
    assign _e_3371 = 37;
    assign _e_3369 = {_e_3370, _e_3371};
    assign _e_3373 = 192;
    assign _e_3374 = 165;
    assign _e_3372 = {_e_3373, _e_3374};
    assign _e_3376 = 192;
    assign _e_3377 = 37;
    assign _e_3375 = {_e_3376, _e_3377};
    assign _e_3379 = 37;
    assign _e_3380 = 0;
    assign _e_3378 = {_e_3379, _e_3380};
    assign _e_3382 = 165;
    assign _e_3383 = 0;
    assign _e_3381 = {_e_3382, _e_3383};
    assign _e_3385 = 165;
    assign _e_3386 = 37;
    assign _e_3384 = {_e_3385, _e_3386};
    assign _e_3388 = 165;
    assign _e_3389 = 165;
    assign _e_3387 = {_e_3388, _e_3389};
    assign _e_3391 = 165;
    assign _e_3392 = 37;
    assign _e_3390 = {_e_3391, _e_3392};
    assign _e_3394 = 37;
    assign _e_3395 = 0;
    assign _e_3393 = {_e_3394, _e_3395};
    assign _e_3397 = 165;
    assign _e_3398 = 0;
    assign _e_3396 = {_e_3397, _e_3398};
    assign _e_3400 = 255;
    assign _e_3401 = 37;
    assign _e_3399 = {_e_3400, _e_3401};
    assign _e_3403 = 255;
    assign _e_3404 = 165;
    assign _e_3402 = {_e_3403, _e_3404};
    assign _e_3406 = 255;
    assign _e_3407 = 37;
    assign _e_3405 = {_e_3406, _e_3407};
    assign _e_3409 = 17;
    assign _e_3410 = 0;
    assign _e_3408 = {_e_3409, _e_3410};
    assign _e_3412 = 145;
    assign _e_3413 = 0;
    assign _e_3411 = {_e_3412, _e_3413};
    assign _e_3415 = 128;
    assign _e_3416 = 61;
    assign _e_3414 = {_e_3415, _e_3416};
    assign _e_3418 = 128;
    assign _e_3419 = 189;
    assign _e_3417 = {_e_3418, _e_3419};
    assign _e_3421 = 128;
    assign _e_3422 = 61;
    assign _e_3420 = {_e_3421, _e_3422};
    assign _e_3424 = 20;
    assign _e_3425 = 0;
    assign _e_3423 = {_e_3424, _e_3425};
    assign _e_3427 = 148;
    assign _e_3428 = 0;
    assign _e_3426 = {_e_3427, _e_3428};
    assign _e_3430 = 145;
    assign _e_3431 = 62;
    assign _e_3429 = {_e_3430, _e_3431};
    assign _e_3433 = 145;
    assign _e_3434 = 190;
    assign _e_3432 = {_e_3433, _e_3434};
    assign _e_3436 = 145;
    assign _e_3437 = 62;
    assign _e_3435 = {_e_3436, _e_3437};
    assign _e_3439 = 20;
    assign _e_3440 = 0;
    assign _e_3438 = {_e_3439, _e_3440};
    assign _e_3442 = 148;
    assign _e_3443 = 0;
    assign _e_3441 = {_e_3442, _e_3443};
    assign _e_3445 = 128;
    assign _e_3446 = 63;
    assign _e_3444 = {_e_3445, _e_3446};
    assign _e_3448 = 128;
    assign _e_3449 = 191;
    assign _e_3447 = {_e_3448, _e_3449};
    assign _e_3451 = 128;
    assign _e_3452 = 63;
    assign _e_3450 = {_e_3451, _e_3452};
    assign _e_3454 = 61;
    assign _e_3455 = 0;
    assign _e_3453 = {_e_3454, _e_3455};
    assign _e_3457 = 189;
    assign _e_3458 = 0;
    assign _e_3456 = {_e_3457, _e_3458};
    assign _e_3460 = 190;
    assign _e_3461 = 20;
    assign _e_3459 = {_e_3460, _e_3461};
    assign _e_3463 = 190;
    assign _e_3464 = 148;
    assign _e_3462 = {_e_3463, _e_3464};
    assign _e_3466 = 190;
    assign _e_3467 = 20;
    assign _e_3465 = {_e_3466, _e_3467};
    assign _e_3469 = 20;
    assign _e_3470 = 0;
    assign _e_3468 = {_e_3469, _e_3470};
    assign _e_3472 = 148;
    assign _e_3473 = 0;
    assign _e_3471 = {_e_3472, _e_3473};
    assign _e_3475 = 148;
    assign _e_3476 = 20;
    assign _e_3474 = {_e_3475, _e_3476};
    assign _e_3478 = 148;
    assign _e_3479 = 148;
    assign _e_3477 = {_e_3478, _e_3479};
    assign _e_3481 = 148;
    assign _e_3482 = 20;
    assign _e_3480 = {_e_3481, _e_3482};
    assign _e_3484 = 20;
    assign _e_3485 = 0;
    assign _e_3483 = {_e_3484, _e_3485};
    assign _e_3487 = 148;
    assign _e_3488 = 0;
    assign _e_3486 = {_e_3487, _e_3488};
    assign _e_3490 = 191;
    assign _e_3491 = 20;
    assign _e_3489 = {_e_3490, _e_3491};
    assign _e_3493 = 191;
    assign _e_3494 = 148;
    assign _e_3492 = {_e_3493, _e_3494};
    assign _e_3496 = 191;
    assign _e_3497 = 20;
    assign _e_3495 = {_e_3496, _e_3497};
    assign _e_3499 = 30;
    assign _e_3500 = 0;
    assign _e_3498 = {_e_3499, _e_3500};
    assign _e_3502 = 158;
    assign _e_3503 = 0;
    assign _e_3501 = {_e_3502, _e_3503};
    assign _e_3505 = 158;
    assign _e_3506 = 10;
    assign _e_3504 = {_e_3505, _e_3506};
    assign _e_3508 = 158;
    assign _e_3509 = 138;
    assign _e_3507 = {_e_3508, _e_3509};
    assign _e_3511 = 158;
    assign _e_3512 = 10;
    assign _e_3510 = {_e_3511, _e_3512};
    assign _e_3514 = 10;
    assign _e_3515 = 1;
    assign _e_3513 = {_e_3514, _e_3515};
    assign _e_3517 = 138;
    assign _e_3518 = 1;
    assign _e_3516 = {_e_3517, _e_3518};
    assign _e_3520 = 138;
    assign _e_3521 = 10;
    assign _e_3519 = {_e_3520, _e_3521};
    assign _e_3523 = 138;
    assign _e_3524 = 138;
    assign _e_3522 = {_e_3523, _e_3524};
    assign _e_3526 = 138;
    assign _e_3527 = 10;
    assign _e_3525 = {_e_3526, _e_3527};
    assign _e_3529 = 31;
    assign _e_3530 = 0;
    assign _e_3528 = {_e_3529, _e_3530};
    assign _e_3532 = 159;
    assign _e_3533 = 0;
    assign _e_3531 = {_e_3532, _e_3533};
    assign _e_3535 = 159;
    assign _e_3536 = 11;
    assign _e_3534 = {_e_3535, _e_3536};
    assign _e_3538 = 159;
    assign _e_3539 = 139;
    assign _e_3537 = {_e_3538, _e_3539};
    assign _e_3541 = 159;
    assign _e_3542 = 11;
    assign _e_3540 = {_e_3541, _e_3542};
    assign _e_3544 = 11;
    assign _e_3545 = 1;
    assign _e_3543 = {_e_3544, _e_3545};
    assign _e_3547 = 139;
    assign _e_3548 = 1;
    assign _e_3546 = {_e_3547, _e_3548};
    assign _e_3550 = 139;
    assign _e_3551 = 11;
    assign _e_3549 = {_e_3550, _e_3551};
    assign _e_3553 = 139;
    assign _e_3554 = 139;
    assign _e_3552 = {_e_3553, _e_3554};
    assign _e_3556 = 139;
    assign _e_3557 = 11;
    assign _e_3555 = {_e_3556, _e_3557};
    assign _e_3559 = 32;
    assign _e_3560 = 0;
    assign _e_3558 = {_e_3559, _e_3560};
    assign _e_3562 = 160;
    assign _e_3563 = 0;
    assign _e_3561 = {_e_3562, _e_3563};
    assign _e_3565 = 160;
    assign _e_3566 = 12;
    assign _e_3564 = {_e_3565, _e_3566};
    assign _e_3568 = 160;
    assign _e_3569 = 140;
    assign _e_3567 = {_e_3568, _e_3569};
    assign _e_3571 = 160;
    assign _e_3572 = 12;
    assign _e_3570 = {_e_3571, _e_3572};
    assign _e_3574 = 12;
    assign _e_3575 = 1;
    assign _e_3573 = {_e_3574, _e_3575};
    assign _e_3577 = 140;
    assign _e_3578 = 1;
    assign _e_3576 = {_e_3577, _e_3578};
    assign _e_3580 = 140;
    assign _e_3581 = 12;
    assign _e_3579 = {_e_3580, _e_3581};
    assign _e_3583 = 140;
    assign _e_3584 = 140;
    assign _e_3582 = {_e_3583, _e_3584};
    assign _e_3586 = 140;
    assign _e_3587 = 12;
    assign _e_3585 = {_e_3586, _e_3587};
    assign _e_3589 = 33;
    assign _e_3590 = 0;
    assign _e_3588 = {_e_3589, _e_3590};
    assign _e_3592 = 161;
    assign _e_3593 = 0;
    assign _e_3591 = {_e_3592, _e_3593};
    assign _e_3595 = 161;
    assign _e_3596 = 13;
    assign _e_3594 = {_e_3595, _e_3596};
    assign _e_3598 = 161;
    assign _e_3599 = 141;
    assign _e_3597 = {_e_3598, _e_3599};
    assign _e_3601 = 161;
    assign _e_3602 = 13;
    assign _e_3600 = {_e_3601, _e_3602};
    assign _e_3604 = 13;
    assign _e_3605 = 1;
    assign _e_3603 = {_e_3604, _e_3605};
    assign _e_3607 = 141;
    assign _e_3608 = 1;
    assign _e_3606 = {_e_3607, _e_3608};
    assign _e_3610 = 141;
    assign _e_3611 = 13;
    assign _e_3609 = {_e_3610, _e_3611};
    assign _e_3613 = 141;
    assign _e_3614 = 141;
    assign _e_3612 = {_e_3613, _e_3614};
    assign _e_3616 = 141;
    assign _e_3617 = 13;
    assign _e_3615 = {_e_3616, _e_3617};
    assign _e_3619 = 34;
    assign _e_3620 = 0;
    assign _e_3618 = {_e_3619, _e_3620};
    assign _e_3622 = 162;
    assign _e_3623 = 0;
    assign _e_3621 = {_e_3622, _e_3623};
    assign _e_3625 = 162;
    assign _e_3626 = 14;
    assign _e_3624 = {_e_3625, _e_3626};
    assign _e_3628 = 162;
    assign _e_3629 = 142;
    assign _e_3627 = {_e_3628, _e_3629};
    assign _e_3631 = 162;
    assign _e_3632 = 14;
    assign _e_3630 = {_e_3631, _e_3632};
    assign _e_3634 = 14;
    assign _e_3635 = 1;
    assign _e_3633 = {_e_3634, _e_3635};
    assign _e_3637 = 142;
    assign _e_3638 = 1;
    assign _e_3636 = {_e_3637, _e_3638};
    assign _e_3640 = 142;
    assign _e_3641 = 14;
    assign _e_3639 = {_e_3640, _e_3641};
    assign _e_3643 = 142;
    assign _e_3644 = 142;
    assign _e_3642 = {_e_3643, _e_3644};
    assign _e_3646 = 142;
    assign _e_3647 = 14;
    assign _e_3645 = {_e_3646, _e_3647};
    assign _e_3649 = 35;
    assign _e_3650 = 0;
    assign _e_3648 = {_e_3649, _e_3650};
    assign _e_3652 = 163;
    assign _e_3653 = 0;
    assign _e_3651 = {_e_3652, _e_3653};
    assign _e_3655 = 163;
    assign _e_3656 = 15;
    assign _e_3654 = {_e_3655, _e_3656};
    assign _e_3658 = 163;
    assign _e_3659 = 143;
    assign _e_3657 = {_e_3658, _e_3659};
    assign _e_3661 = 163;
    assign _e_3662 = 15;
    assign _e_3660 = {_e_3661, _e_3662};
    assign _e_3664 = 15;
    assign _e_3665 = 1;
    assign _e_3663 = {_e_3664, _e_3665};
    assign _e_3667 = 143;
    assign _e_3668 = 1;
    assign _e_3666 = {_e_3667, _e_3668};
    assign _e_3670 = 143;
    assign _e_3671 = 15;
    assign _e_3669 = {_e_3670, _e_3671};
    assign _e_3673 = 143;
    assign _e_3674 = 143;
    assign _e_3672 = {_e_3673, _e_3674};
    assign _e_3676 = 143;
    assign _e_3677 = 15;
    assign _e_3675 = {_e_3676, _e_3677};
    assign _e_3679 = 36;
    assign _e_3680 = 0;
    assign _e_3678 = {_e_3679, _e_3680};
    assign _e_3682 = 164;
    assign _e_3683 = 0;
    assign _e_3681 = {_e_3682, _e_3683};
    assign _e_3685 = 164;
    assign _e_3686 = 16;
    assign _e_3684 = {_e_3685, _e_3686};
    assign _e_3688 = 164;
    assign _e_3689 = 144;
    assign _e_3687 = {_e_3688, _e_3689};
    assign _e_3691 = 164;
    assign _e_3692 = 16;
    assign _e_3690 = {_e_3691, _e_3692};
    assign _e_3694 = 16;
    assign _e_3695 = 1;
    assign _e_3693 = {_e_3694, _e_3695};
    assign _e_3697 = 144;
    assign _e_3698 = 1;
    assign _e_3696 = {_e_3697, _e_3698};
    assign _e_3700 = 144;
    assign _e_3701 = 16;
    assign _e_3699 = {_e_3700, _e_3701};
    assign _e_3703 = 144;
    assign _e_3704 = 144;
    assign _e_3702 = {_e_3703, _e_3704};
    assign _e_3706 = 144;
    assign _e_3707 = 16;
    assign _e_3705 = {_e_3706, _e_3707};
    assign _e_3709 = 37;
    assign _e_3710 = 0;
    assign _e_3708 = {_e_3709, _e_3710};
    assign _e_3712 = 165;
    assign _e_3713 = 0;
    assign _e_3711 = {_e_3712, _e_3713};
    assign _e_3715 = 165;
    assign _e_3716 = 17;
    assign _e_3714 = {_e_3715, _e_3716};
    assign _e_3718 = 165;
    assign _e_3719 = 145;
    assign _e_3717 = {_e_3718, _e_3719};
    assign _e_3721 = 165;
    assign _e_3722 = 17;
    assign _e_3720 = {_e_3721, _e_3722};
    assign _e_3724 = 17;
    assign _e_3725 = 1;
    assign _e_3723 = {_e_3724, _e_3725};
    assign _e_3727 = 145;
    assign _e_3728 = 1;
    assign _e_3726 = {_e_3727, _e_3728};
    assign _e_3730 = 145;
    assign _e_3731 = 17;
    assign _e_3729 = {_e_3730, _e_3731};
    assign _e_3733 = 145;
    assign _e_3734 = 145;
    assign _e_3732 = {_e_3733, _e_3734};
    assign _e_3736 = 145;
    assign _e_3737 = 17;
    assign _e_3735 = {_e_3736, _e_3737};
    assign _e_362 = {_e_3735, _e_3732, _e_3729, _e_3726, _e_3723, _e_3720, _e_3717, _e_3714, _e_3711, _e_3708, _e_3705, _e_3702, _e_3699, _e_3696, _e_3693, _e_3690, _e_3687, _e_3684, _e_3681, _e_3678, _e_3675, _e_3672, _e_3669, _e_3666, _e_3663, _e_3660, _e_3657, _e_3654, _e_3651, _e_3648, _e_3645, _e_3642, _e_3639, _e_3636, _e_3633, _e_3630, _e_3627, _e_3624, _e_3621, _e_3618, _e_3615, _e_3612, _e_3609, _e_3606, _e_3603, _e_3600, _e_3597, _e_3594, _e_3591, _e_3588, _e_3585, _e_3582, _e_3579, _e_3576, _e_3573, _e_3570, _e_3567, _e_3564, _e_3561, _e_3558, _e_3555, _e_3552, _e_3549, _e_3546, _e_3543, _e_3540, _e_3537, _e_3534, _e_3531, _e_3528, _e_3525, _e_3522, _e_3519, _e_3516, _e_3513, _e_3510, _e_3507, _e_3504, _e_3501, _e_3498, _e_3495, _e_3492, _e_3489, _e_3486, _e_3483, _e_3480, _e_3477, _e_3474, _e_3471, _e_3468, _e_3465, _e_3462, _e_3459, _e_3456, _e_3453, _e_3450, _e_3447, _e_3444, _e_3441, _e_3438, _e_3435, _e_3432, _e_3429, _e_3426, _e_3423, _e_3420, _e_3417, _e_3414, _e_3411, _e_3408, _e_3405, _e_3402, _e_3399, _e_3396, _e_3393, _e_3390, _e_3387, _e_3384, _e_3381, _e_3378, _e_3375, _e_3372, _e_3369, _e_3366, _e_3363, _e_3360, _e_3357, _e_3354, _e_3351, _e_3348, _e_3345, _e_3342, _e_3339, _e_3336, _e_3333, _e_3330, _e_3327, _e_3324, _e_3321, _e_3318, _e_3315, _e_3312, _e_3309, _e_3306, _e_3303, _e_3300, _e_3297, _e_3294, _e_3291, _e_3288, _e_3285, _e_3282, _e_3279, _e_3276, _e_3273, _e_3270, _e_3267, _e_3264, _e_3261, _e_3258, _e_3255, _e_3252, _e_3249, _e_3246, _e_3243, _e_3240, _e_3237, _e_3234, _e_3231, _e_3228, _e_3225, _e_3222, _e_3219, _e_3216, _e_3213, _e_3210, _e_3207, _e_3204, _e_3201, _e_3198, _e_3195, _e_3192, _e_3189, _e_3186, _e_3183, _e_3180, _e_3177, _e_3174, _e_3171, _e_3168, _e_3165, _e_3162, _e_3159, _e_3156, _e_3153, _e_3150, _e_3147, _e_3144, _e_3141, _e_3138, _e_3135, _e_3132, _e_3129, _e_3126, _e_3123, _e_3120, _e_3117, _e_3114, _e_3111, _e_3108, _e_3105, _e_3102, _e_3099, _e_3096, _e_3093, _e_3090, _e_3087, _e_3084, _e_3081, _e_3078, _e_3075, _e_3072, _e_3069, _e_3066, _e_3063, _e_3060, _e_3057, _e_3054, _e_3051, _e_3048, _e_3045, _e_3042, _e_3039, _e_3036, _e_3033, _e_3030, _e_3027, _e_3024, _e_3021, _e_3018, _e_3015, _e_3012, _e_3009, _e_3006, _e_3003, _e_3000, _e_2997, _e_2994, _e_2991, _e_2988, _e_2985, _e_2982, _e_2979, _e_2976, _e_2973, _e_2970, _e_2967, _e_2964, _e_2961, _e_2958, _e_2955, _e_2952, _e_2949, _e_2946, _e_2943, _e_2940, _e_2937, _e_2934, _e_2931, _e_2928, _e_2925, _e_2922, _e_2919, _e_2916, _e_2913, _e_2910, _e_2907, _e_2904, _e_2901, _e_2898, _e_2895, _e_2892, _e_2889, _e_2886, _e_2883, _e_2880, _e_2877, _e_2874, _e_2871, _e_2868, _e_2865, _e_2862, _e_2859, _e_2856, _e_2853, _e_2850, _e_2847, _e_2844, _e_2841, _e_2838, _e_2835, _e_2832, _e_2829, _e_2826, _e_2823, _e_2820, _e_2817, _e_2814, _e_2811, _e_2808, _e_2805, _e_2802, _e_2799, _e_2796, _e_2793, _e_2790, _e_2787, _e_2784, _e_2781, _e_2778, _e_2775, _e_2772, _e_2769, _e_2766, _e_2763, _e_2760, _e_2757, _e_2754, _e_2751, _e_2748, _e_2745, _e_2742, _e_2739, _e_2736, _e_2733, _e_2730, _e_2727, _e_2724, _e_2721, _e_2718, _e_2715, _e_2712, _e_2709, _e_2706, _e_2703, _e_2700, _e_2697, _e_2694, _e_2691, _e_2688, _e_2685, _e_2682, _e_2679, _e_2676, _e_2673, _e_2670, _e_2667, _e_2664, _e_2661, _e_2658, _e_2655, _e_2652, _e_2649, _e_2646, _e_2643, _e_2640, _e_2637, _e_2634, _e_2631, _e_2628, _e_2625, _e_2622, _e_2619, _e_2616, _e_2613, _e_2610, _e_2607, _e_2604, _e_2601, _e_2598, _e_2595, _e_2592, _e_2589, _e_2586, _e_2583, _e_2580, _e_2577, _e_2574, _e_2571, _e_2568, _e_2565, _e_2562, _e_2559, _e_2556, _e_2553, _e_2550, _e_2547, _e_2544, _e_2541, _e_2538, _e_2535, _e_2532, _e_2529, _e_2526, _e_2523, _e_2520, _e_2517, _e_2514, _e_2511, _e_2508, _e_2505, _e_2502, _e_2499, _e_2496, _e_2493, _e_2490, _e_2487, _e_2484, _e_2481, _e_2478, _e_2475, _e_2472, _e_2469, _e_2466, _e_2463, _e_2460, _e_2457, _e_2454, _e_2451, _e_2448, _e_2445, _e_2442, _e_2439, _e_2436, _e_2433, _e_2430, _e_2427, _e_2424, _e_2421, _e_2418, _e_2415, _e_2412, _e_2409, _e_2406, _e_2403, _e_2400, _e_2397, _e_2394, _e_2391, _e_2388, _e_2385, _e_2382, _e_2379, _e_2376, _e_2373, _e_2370, _e_2367, _e_2364, _e_2361, _e_2358, _e_2355, _e_2352, _e_2349, _e_2346, _e_2343, _e_2340, _e_2337, _e_2334, _e_2331, _e_2328, _e_2325, _e_2322, _e_2319, _e_2316, _e_2313, _e_2310, _e_2307, _e_2304, _e_2301, _e_2298, _e_2295, _e_2292, _e_2289, _e_2286, _e_2283, _e_2280, _e_2277, _e_2274, _e_2271, _e_2268, _e_2265, _e_2262, _e_2259, _e_2256, _e_2253, _e_2250, _e_2247, _e_2244, _e_2241, _e_2238, _e_2235, _e_2232, _e_2229, _e_2226, _e_2223, _e_2220, _e_2217, _e_2214, _e_2211, _e_2208, _e_2205, _e_2202, _e_2199, _e_2196, _e_2193, _e_2190, _e_2187, _e_2184, _e_2181, _e_2178, _e_2175, _e_2172, _e_2169, _e_2166, _e_2163, _e_2160, _e_2157, _e_2154, _e_2151, _e_2148, _e_2145, _e_2142, _e_2139, _e_2136, _e_2133, _e_2130, _e_2127, _e_2124, _e_2121, _e_2118, _e_2115, _e_2112, _e_2109, _e_2106, _e_2103, _e_2100, _e_2097, _e_2094, _e_2091, _e_2088, _e_2085, _e_2082, _e_2079, _e_2076, _e_2073, _e_2070, _e_2067, _e_2064, _e_2061, _e_2058, _e_2055, _e_2052, _e_2049, _e_2046, _e_2043, _e_2040, _e_2037, _e_2034, _e_2031, _e_2028, _e_2025, _e_2022, _e_2019, _e_2016, _e_2013, _e_2010, _e_2007, _e_2004, _e_2001, _e_1998, _e_1995, _e_1992, _e_1989, _e_1986, _e_1983, _e_1980, _e_1977, _e_1974, _e_1971, _e_1968, _e_1965, _e_1962, _e_1959, _e_1956, _e_1953, _e_1950, _e_1947, _e_1944, _e_1941, _e_1938, _e_1935, _e_1932, _e_1929, _e_1926, _e_1923, _e_1920, _e_1917, _e_1914, _e_1911, _e_1908, _e_1905, _e_1902, _e_1899, _e_1896, _e_1893, _e_1890, _e_1887, _e_1884, _e_1881, _e_1878, _e_1875, _e_1872, _e_1869, _e_1866, _e_1863, _e_1860, _e_1857, _e_1854, _e_1851, _e_1848, _e_1845, _e_1842, _e_1839, _e_1836, _e_1833, _e_1830, _e_1827, _e_1824, _e_1821, _e_1818, _e_1815, _e_1812, _e_1809, _e_1806, _e_1803, _e_1800, _e_1797, _e_1794, _e_1791, _e_1788, _e_1785, _e_1782, _e_1779, _e_1776, _e_1773, _e_1770, _e_1767, _e_1764, _e_1761, _e_1758, _e_1755, _e_1752, _e_1749, _e_1746, _e_1743, _e_1740, _e_1737, _e_1734, _e_1731, _e_1728, _e_1725, _e_1722, _e_1719, _e_1716, _e_1713, _e_1710, _e_1707, _e_1704, _e_1701, _e_1698, _e_1695, _e_1692, _e_1689, _e_1686, _e_1683, _e_1680, _e_1677, _e_1674, _e_1671, _e_1668, _e_1665, _e_1662, _e_1659, _e_1656, _e_1653, _e_1650, _e_1647, _e_1644, _e_1641, _e_1638, _e_1635, _e_1632, _e_1629, _e_1626, _e_1623, _e_1620, _e_1617, _e_1614, _e_1611, _e_1608, _e_1605, _e_1602, _e_1599, _e_1596, _e_1593, _e_1590, _e_1587, _e_1584, _e_1581, _e_1578, _e_1575, _e_1572, _e_1569, _e_1566, _e_1563, _e_1560, _e_1557, _e_1554, _e_1551, _e_1548, _e_1545, _e_1542, _e_1539, _e_1536, _e_1533, _e_1530, _e_1527, _e_1524, _e_1521, _e_1518, _e_1515, _e_1512, _e_1509, _e_1506, _e_1503, _e_1500, _e_1497, _e_1494, _e_1491, _e_1488, _e_1485, _e_1482, _e_1479, _e_1476, _e_1473, _e_1470, _e_1467, _e_1464, _e_1461, _e_1458, _e_1455, _e_1452, _e_1449, _e_1446, _e_1443, _e_1440, _e_1437, _e_1434, _e_1431, _e_1428, _e_1425, _e_1422, _e_1419, _e_1416, _e_1413, _e_1410, _e_1407, _e_1404, _e_1401, _e_1398, _e_1395, _e_1392, _e_1389, _e_1386, _e_1383, _e_1380, _e_1377, _e_1374, _e_1371, _e_1368, _e_1365, _e_1362, _e_1359, _e_1356, _e_1353, _e_1350, _e_1347, _e_1344, _e_1341, _e_1338, _e_1335, _e_1332, _e_1329, _e_1326, _e_1323, _e_1320, _e_1317, _e_1314, _e_1311, _e_1308, _e_1305, _e_1302, _e_1299, _e_1296, _e_1293, _e_1290, _e_1287, _e_1284, _e_1281, _e_1278, _e_1275, _e_1272, _e_1269, _e_1266, _e_1263, _e_1260, _e_1257, _e_1254, _e_1251, _e_1248, _e_1245, _e_1242, _e_1239, _e_1236, _e_1233, _e_1230, _e_1227, _e_1224, _e_1221, _e_1218, _e_1215, _e_1212, _e_1209, _e_1206, _e_1203, _e_1200, _e_1197, _e_1194, _e_1191, _e_1188, _e_1185, _e_1182, _e_1179, _e_1176, _e_1173, _e_1170, _e_1167, _e_1164, _e_1161, _e_1158, _e_1155, _e_1152, _e_1149, _e_1146, _e_1143, _e_1140, _e_1137, _e_1134, _e_1131, _e_1128, _e_1125, _e_1122, _e_1119, _e_1116, _e_1113, _e_1110, _e_1107, _e_1104, _e_1101, _e_1098, _e_1095, _e_1092, _e_1089, _e_1086, _e_1083, _e_1080, _e_1077, _e_1074, _e_1071, _e_1068, _e_1065, _e_1062, _e_1059, _e_1056, _e_1053, _e_1050, _e_1047, _e_1044, _e_1041, _e_1038, _e_1035, _e_1032, _e_1029, _e_1026, _e_1023, _e_1020, _e_1017, _e_1014, _e_1011, _e_1008, _e_1005, _e_1002, _e_999, _e_996, _e_993, _e_990, _e_987, _e_984, _e_981, _e_978, _e_975, _e_972, _e_969, _e_966, _e_963, _e_960, _e_957, _e_954, _e_951, _e_948, _e_945, _e_942, _e_939, _e_936, _e_933, _e_930, _e_927, _e_924, _e_921, _e_918, _e_915, _e_912, _e_909, _e_906, _e_903, _e_900, _e_897, _e_894, _e_891, _e_888, _e_885, _e_882, _e_879, _e_876, _e_873, _e_870, _e_867, _e_864, _e_861, _e_858, _e_855, _e_852, _e_849, _e_846, _e_843, _e_840, _e_837, _e_834, _e_831, _e_828, _e_825, _e_822, _e_819, _e_816, _e_813, _e_810, _e_807, _e_804, _e_801, _e_798, _e_795, _e_792, _e_789, _e_786, _e_783, _e_780, _e_777, _e_774, _e_771, _e_768, _e_765, _e_762, _e_759, _e_756, _e_753, _e_750, _e_747, _e_744, _e_741, _e_738, _e_735, _e_732, _e_729, _e_726, _e_723, _e_720, _e_717, _e_714, _e_711, _e_708, _e_705, _e_702, _e_699, _e_696, _e_693, _e_690, _e_687, _e_684, _e_681, _e_678, _e_675, _e_672, _e_669, _e_666, _e_663, _e_660, _e_657, _e_654, _e_651, _e_648, _e_645, _e_642, _e_639, _e_636, _e_633, _e_630, _e_627, _e_624, _e_621, _e_618, _e_615, _e_612, _e_609, _e_606, _e_603, _e_600, _e_597, _e_594, _e_591, _e_588, _e_585, _e_582, _e_579, _e_576, _e_573, _e_570, _e_567, _e_564, _e_561, _e_558, _e_555, _e_552, _e_549, _e_546, _e_543, _e_540, _e_537, _e_534, _e_531, _e_528, _e_525, _e_522, _e_519, _e_516, _e_513, _e_510, _e_507, _e_504, _e_501, _e_498, _e_495, _e_492, _e_489, _e_486, _e_483, _e_480, _e_477, _e_474, _e_471, _e_468, _e_465, _e_462, _e_459, _e_456, _e_453, _e_450, _e_447, _e_444, _e_441, _e_438, _e_435, _e_432, _e_429, _e_426, _e_423, _e_420, _e_417, _e_414, _e_411, _e_408, _e_405, _e_402, _e_399, _e_396, _e_393, _e_390, _e_387, _e_384, _e_381, _e_378, _e_375, _e_372, _e_369, _e_366, _e_363};
    initial begin
        \commands [0] = 'b0000000000000000;
        \commands [1] = 'b1000000000000000;
        \commands [2] = 'b1000000000010100;
        \commands [3] = 'b1000000010010100;
        \commands [4] = 'b1000000000010100;
        \commands [5] = 'b0000101000000000;
        \commands [6] = 'b1000101000000000;
        \commands [7] = 'b1000101000110010;
        \commands [8] = 'b1000101010110010;
        \commands [9] = 'b1000101000110010;
        \commands [10] = 'b0000000000000000;
        \commands [11] = 'b1000000000000000;
        \commands [12] = 'b1000000000110011;
        \commands [13] = 'b1000000010110011;
        \commands [14] = 'b1000000000110011;
        \commands [15] = 'b0001010000000000;
        \commands [16] = 'b1001010000000000;
        \commands [17] = 'b1001010000110100;
        \commands [18] = 'b1001010010110100;
        \commands [19] = 'b1001010000110100;
        \commands [20] = 'b0001010000000000;
        \commands [21] = 'b1001010000000000;
        \commands [22] = 'b1011001000111101;
        \commands [23] = 'b1011001010111101;
        \commands [24] = 'b1011001000111101;
        \commands [25] = 'b0011110100000000;
        \commands [26] = 'b1011110100000000;
        \commands [27] = 'b1011110100111101;
        \commands [28] = 'b1011110110111101;
        \commands [29] = 'b1011110100111101;
        \commands [30] = 'b0011110100000000;
        \commands [31] = 'b1011110100000000;
        \commands [32] = 'b1011001100111101;
        \commands [33] = 'b1011001110111101;
        \commands [34] = 'b1011001100111101;
        \commands [35] = 'b0011010000000000;
        \commands [36] = 'b1011010000000000;
        \commands [37] = 'b1011001000111110;
        \commands [38] = 'b1011001010111110;
        \commands [39] = 'b1011001000111110;
        \commands [40] = 'b0011111000000000;
        \commands [41] = 'b1011111000000000;
        \commands [42] = 'b1011111000111110;
        \commands [43] = 'b1011111010111110;
        \commands [44] = 'b1011111000111110;
        \commands [45] = 'b0011111000000000;
        \commands [46] = 'b1011111000000000;
        \commands [47] = 'b1000000000111110;
        \commands [48] = 'b1000000010111110;
        \commands [49] = 'b1000000000111110;
        \commands [50] = 'b0001010000000000;
        \commands [51] = 'b1001010000000000;
        \commands [52] = 'b1000101000111111;
        \commands [53] = 'b1000101010111111;
        \commands [54] = 'b1000101000111111;
        \commands [55] = 'b0011111100000000;
        \commands [56] = 'b1011111100000000;
        \commands [57] = 'b1011111100111111;
        \commands [58] = 'b1011111110111111;
        \commands [59] = 'b1011111100111111;
        \commands [60] = 'b0011111100000000;
        \commands [61] = 'b1011111100000000;
        \commands [62] = 'b1000000000111111;
        \commands [63] = 'b1000000010111111;
        \commands [64] = 'b1000000000111111;
        \commands [65] = 'b0011010000000000;
        \commands [66] = 'b1011010000000000;
        \commands [67] = 'b1000101001000000;
        \commands [68] = 'b1000101011000000;
        \commands [69] = 'b1000101001000000;
        \commands [70] = 'b0100000000000000;
        \commands [71] = 'b1100000000000000;
        \commands [72] = 'b1100000001000000;
        \commands [73] = 'b1100000011000000;
        \commands [74] = 'b1100000001000000;
        \commands [75] = 'b0100000000000000;
        \commands [76] = 'b1100000000000000;
        \commands [77] = 'b1011001101000000;
        \commands [78] = 'b1011001111000000;
        \commands [79] = 'b1011001101000000;
        \commands [80] = 'b0011110100000000;
        \commands [81] = 'b1011110100000000;
        \commands [82] = 'b1011111001111111;
        \commands [83] = 'b1011111011111111;
        \commands [84] = 'b1011111001111111;
        \commands [85] = 'b0111111100000000;
        \commands [86] = 'b1111111100000000;
        \commands [87] = 'b1111111101111111;
        \commands [88] = 'b1111111111111111;
        \commands [89] = 'b1111111101111111;
        \commands [90] = 'b0011111100000000;
        \commands [91] = 'b1011111100000000;
        \commands [92] = 'b1100000000011110;
        \commands [93] = 'b1100000010011110;
        \commands [94] = 'b1100000000011110;
        \commands [95] = 'b0001111000000000;
        \commands [96] = 'b1001111000000000;
        \commands [97] = 'b1001111000011110;
        \commands [98] = 'b1001111010011110;
        \commands [99] = 'b1001111000011110;
        \commands [100] = 'b0001111000000000;
        \commands [101] = 'b1001111000000000;
        \commands [102] = 'b1111111100011110;
        \commands [103] = 'b1111111110011110;
        \commands [104] = 'b1111111100011110;
        \commands [105] = 'b0000101000000000;
        \commands [106] = 'b1000101000000000;
        \commands [107] = 'b1000000000111101;
        \commands [108] = 'b1000000010111101;
        \commands [109] = 'b1000000000111101;
        \commands [110] = 'b0001010000000000;
        \commands [111] = 'b1001010000000000;
        \commands [112] = 'b1000101000111110;
        \commands [113] = 'b1000101010111110;
        \commands [114] = 'b1000101000111110;
        \commands [115] = 'b0001010000000000;
        \commands [116] = 'b1001010000000000;
        \commands [117] = 'b1000000000111111;
        \commands [118] = 'b1000000010111111;
        \commands [119] = 'b1000000000111111;
        \commands [120] = 'b0011110100000000;
        \commands [121] = 'b1011110100000000;
        \commands [122] = 'b1011111000010100;
        \commands [123] = 'b1011111010010100;
        \commands [124] = 'b1011111000010100;
        \commands [125] = 'b0001010000000000;
        \commands [126] = 'b1001010000000000;
        \commands [127] = 'b1001010000010100;
        \commands [128] = 'b1001010010010100;
        \commands [129] = 'b1001010000010100;
        \commands [130] = 'b0001010000000000;
        \commands [131] = 'b1001010000000000;
        \commands [132] = 'b1011111100010100;
        \commands [133] = 'b1011111110010100;
        \commands [134] = 'b1011111100010100;
        \commands [135] = 'b0000101100000000;
        \commands [136] = 'b1000101100000000;
        \commands [137] = 'b1000101100110010;
        \commands [138] = 'b1000101110110010;
        \commands [139] = 'b1000101100110010;
        \commands [140] = 'b0000000000000000;
        \commands [141] = 'b1000000000000000;
        \commands [142] = 'b1000000000110011;
        \commands [143] = 'b1000000010110011;
        \commands [144] = 'b1000000000110011;
        \commands [145] = 'b0001010000000000;
        \commands [146] = 'b1001010000000000;
        \commands [147] = 'b1001010000110100;
        \commands [148] = 'b1001010010110100;
        \commands [149] = 'b1001010000110100;
        \commands [150] = 'b0001010000000000;
        \commands [151] = 'b1001010000000000;
        \commands [152] = 'b1011001000111101;
        \commands [153] = 'b1011001010111101;
        \commands [154] = 'b1011001000111101;
        \commands [155] = 'b0011110100000000;
        \commands [156] = 'b1011110100000000;
        \commands [157] = 'b1011110100111101;
        \commands [158] = 'b1011110110111101;
        \commands [159] = 'b1011110100111101;
        \commands [160] = 'b0011110100000000;
        \commands [161] = 'b1011110100000000;
        \commands [162] = 'b1011001100111101;
        \commands [163] = 'b1011001110111101;
        \commands [164] = 'b1011001100111101;
        \commands [165] = 'b0011010000000000;
        \commands [166] = 'b1011010000000000;
        \commands [167] = 'b1011001000111110;
        \commands [168] = 'b1011001010111110;
        \commands [169] = 'b1011001000111110;
        \commands [170] = 'b0011111000000000;
        \commands [171] = 'b1011111000000000;
        \commands [172] = 'b1011111000111110;
        \commands [173] = 'b1011111010111110;
        \commands [174] = 'b1011111000111110;
        \commands [175] = 'b0011111000000000;
        \commands [176] = 'b1011111000000000;
        \commands [177] = 'b1000000000111110;
        \commands [178] = 'b1000000010111110;
        \commands [179] = 'b1000000000111110;
        \commands [180] = 'b0001010000000000;
        \commands [181] = 'b1001010000000000;
        \commands [182] = 'b1000101100111111;
        \commands [183] = 'b1000101110111111;
        \commands [184] = 'b1000101100111111;
        \commands [185] = 'b0011111100000000;
        \commands [186] = 'b1011111100000000;
        \commands [187] = 'b1011111100111111;
        \commands [188] = 'b1011111110111111;
        \commands [189] = 'b1011111100111111;
        \commands [190] = 'b0011111100000000;
        \commands [191] = 'b1011111100000000;
        \commands [192] = 'b1000000000111111;
        \commands [193] = 'b1000000010111111;
        \commands [194] = 'b1000000000111111;
        \commands [195] = 'b0011010000000000;
        \commands [196] = 'b1011010000000000;
        \commands [197] = 'b1000101101000000;
        \commands [198] = 'b1000101111000000;
        \commands [199] = 'b1000101101000000;
        \commands [200] = 'b0100000000000000;
        \commands [201] = 'b1100000000000000;
        \commands [202] = 'b1100000001000000;
        \commands [203] = 'b1100000011000000;
        \commands [204] = 'b1100000001000000;
        \commands [205] = 'b0100000000000000;
        \commands [206] = 'b1100000000000000;
        \commands [207] = 'b1011001101000000;
        \commands [208] = 'b1011001111000000;
        \commands [209] = 'b1011001101000000;
        \commands [210] = 'b0011110100000000;
        \commands [211] = 'b1011110100000000;
        \commands [212] = 'b1011111001111111;
        \commands [213] = 'b1011111011111111;
        \commands [214] = 'b1011111001111111;
        \commands [215] = 'b0111111100000000;
        \commands [216] = 'b1111111100000000;
        \commands [217] = 'b1111111101111111;
        \commands [218] = 'b1111111111111111;
        \commands [219] = 'b1111111101111111;
        \commands [220] = 'b0011111100000000;
        \commands [221] = 'b1011111100000000;
        \commands [222] = 'b1100000000011111;
        \commands [223] = 'b1100000010011111;
        \commands [224] = 'b1100000000011111;
        \commands [225] = 'b0001111100000000;
        \commands [226] = 'b1001111100000000;
        \commands [227] = 'b1001111100011111;
        \commands [228] = 'b1001111110011111;
        \commands [229] = 'b1001111100011111;
        \commands [230] = 'b0001111100000000;
        \commands [231] = 'b1001111100000000;
        \commands [232] = 'b1111111100011111;
        \commands [233] = 'b1111111110011111;
        \commands [234] = 'b1111111100011111;
        \commands [235] = 'b0000101100000000;
        \commands [236] = 'b1000101100000000;
        \commands [237] = 'b1000000000111101;
        \commands [238] = 'b1000000010111101;
        \commands [239] = 'b1000000000111101;
        \commands [240] = 'b0001010000000000;
        \commands [241] = 'b1001010000000000;
        \commands [242] = 'b1000101100111110;
        \commands [243] = 'b1000101110111110;
        \commands [244] = 'b1000101100111110;
        \commands [245] = 'b0001010000000000;
        \commands [246] = 'b1001010000000000;
        \commands [247] = 'b1000000000111111;
        \commands [248] = 'b1000000010111111;
        \commands [249] = 'b1000000000111111;
        \commands [250] = 'b0011110100000000;
        \commands [251] = 'b1011110100000000;
        \commands [252] = 'b1011111000010100;
        \commands [253] = 'b1011111010010100;
        \commands [254] = 'b1011111000010100;
        \commands [255] = 'b0001010000000000;
        \commands [256] = 'b1001010000000000;
        \commands [257] = 'b1001010000010100;
        \commands [258] = 'b1001010010010100;
        \commands [259] = 'b1001010000010100;
        \commands [260] = 'b0001010000000000;
        \commands [261] = 'b1001010000000000;
        \commands [262] = 'b1011111100010100;
        \commands [263] = 'b1011111110010100;
        \commands [264] = 'b1011111100010100;
        \commands [265] = 'b0000110000000000;
        \commands [266] = 'b1000110000000000;
        \commands [267] = 'b1000110000110010;
        \commands [268] = 'b1000110010110010;
        \commands [269] = 'b1000110000110010;
        \commands [270] = 'b0000000000000000;
        \commands [271] = 'b1000000000000000;
        \commands [272] = 'b1000000000110011;
        \commands [273] = 'b1000000010110011;
        \commands [274] = 'b1000000000110011;
        \commands [275] = 'b0001010000000000;
        \commands [276] = 'b1001010000000000;
        \commands [277] = 'b1001010000110100;
        \commands [278] = 'b1001010010110100;
        \commands [279] = 'b1001010000110100;
        \commands [280] = 'b0001010000000000;
        \commands [281] = 'b1001010000000000;
        \commands [282] = 'b1011001000111101;
        \commands [283] = 'b1011001010111101;
        \commands [284] = 'b1011001000111101;
        \commands [285] = 'b0011110100000000;
        \commands [286] = 'b1011110100000000;
        \commands [287] = 'b1011110100111101;
        \commands [288] = 'b1011110110111101;
        \commands [289] = 'b1011110100111101;
        \commands [290] = 'b0011110100000000;
        \commands [291] = 'b1011110100000000;
        \commands [292] = 'b1011001100111101;
        \commands [293] = 'b1011001110111101;
        \commands [294] = 'b1011001100111101;
        \commands [295] = 'b0011010000000000;
        \commands [296] = 'b1011010000000000;
        \commands [297] = 'b1011001000111110;
        \commands [298] = 'b1011001010111110;
        \commands [299] = 'b1011001000111110;
        \commands [300] = 'b0011111000000000;
        \commands [301] = 'b1011111000000000;
        \commands [302] = 'b1011111000111110;
        \commands [303] = 'b1011111010111110;
        \commands [304] = 'b1011111000111110;
        \commands [305] = 'b0011111000000000;
        \commands [306] = 'b1011111000000000;
        \commands [307] = 'b1000000000111110;
        \commands [308] = 'b1000000010111110;
        \commands [309] = 'b1000000000111110;
        \commands [310] = 'b0001010000000000;
        \commands [311] = 'b1001010000000000;
        \commands [312] = 'b1000110000111111;
        \commands [313] = 'b1000110010111111;
        \commands [314] = 'b1000110000111111;
        \commands [315] = 'b0011111100000000;
        \commands [316] = 'b1011111100000000;
        \commands [317] = 'b1011111100111111;
        \commands [318] = 'b1011111110111111;
        \commands [319] = 'b1011111100111111;
        \commands [320] = 'b0011111100000000;
        \commands [321] = 'b1011111100000000;
        \commands [322] = 'b1000000000111111;
        \commands [323] = 'b1000000010111111;
        \commands [324] = 'b1000000000111111;
        \commands [325] = 'b0011010000000000;
        \commands [326] = 'b1011010000000000;
        \commands [327] = 'b1000110001000000;
        \commands [328] = 'b1000110011000000;
        \commands [329] = 'b1000110001000000;
        \commands [330] = 'b0100000000000000;
        \commands [331] = 'b1100000000000000;
        \commands [332] = 'b1100000001000000;
        \commands [333] = 'b1100000011000000;
        \commands [334] = 'b1100000001000000;
        \commands [335] = 'b0100000000000000;
        \commands [336] = 'b1100000000000000;
        \commands [337] = 'b1011001101000000;
        \commands [338] = 'b1011001111000000;
        \commands [339] = 'b1011001101000000;
        \commands [340] = 'b0011110100000000;
        \commands [341] = 'b1011110100000000;
        \commands [342] = 'b1011111001111111;
        \commands [343] = 'b1011111011111111;
        \commands [344] = 'b1011111001111111;
        \commands [345] = 'b0111111100000000;
        \commands [346] = 'b1111111100000000;
        \commands [347] = 'b1111111101111111;
        \commands [348] = 'b1111111111111111;
        \commands [349] = 'b1111111101111111;
        \commands [350] = 'b0011111100000000;
        \commands [351] = 'b1011111100000000;
        \commands [352] = 'b1100000000100000;
        \commands [353] = 'b1100000010100000;
        \commands [354] = 'b1100000000100000;
        \commands [355] = 'b0010000000000000;
        \commands [356] = 'b1010000000000000;
        \commands [357] = 'b1010000000100000;
        \commands [358] = 'b1010000010100000;
        \commands [359] = 'b1010000000100000;
        \commands [360] = 'b0010000000000000;
        \commands [361] = 'b1010000000000000;
        \commands [362] = 'b1111111100100000;
        \commands [363] = 'b1111111110100000;
        \commands [364] = 'b1111111100100000;
        \commands [365] = 'b0000110000000000;
        \commands [366] = 'b1000110000000000;
        \commands [367] = 'b1000000000111101;
        \commands [368] = 'b1000000010111101;
        \commands [369] = 'b1000000000111101;
        \commands [370] = 'b0001010000000000;
        \commands [371] = 'b1001010000000000;
        \commands [372] = 'b1000110000111110;
        \commands [373] = 'b1000110010111110;
        \commands [374] = 'b1000110000111110;
        \commands [375] = 'b0001010000000000;
        \commands [376] = 'b1001010000000000;
        \commands [377] = 'b1000000000111111;
        \commands [378] = 'b1000000010111111;
        \commands [379] = 'b1000000000111111;
        \commands [380] = 'b0011110100000000;
        \commands [381] = 'b1011110100000000;
        \commands [382] = 'b1011111000010100;
        \commands [383] = 'b1011111010010100;
        \commands [384] = 'b1011111000010100;
        \commands [385] = 'b0001010000000000;
        \commands [386] = 'b1001010000000000;
        \commands [387] = 'b1001010000010100;
        \commands [388] = 'b1001010010010100;
        \commands [389] = 'b1001010000010100;
        \commands [390] = 'b0001010000000000;
        \commands [391] = 'b1001010000000000;
        \commands [392] = 'b1011111100010100;
        \commands [393] = 'b1011111110010100;
        \commands [394] = 'b1011111100010100;
        \commands [395] = 'b0000110100000000;
        \commands [396] = 'b1000110100000000;
        \commands [397] = 'b1000110100110010;
        \commands [398] = 'b1000110110110010;
        \commands [399] = 'b1000110100110010;
        \commands [400] = 'b0000000000000000;
        \commands [401] = 'b1000000000000000;
        \commands [402] = 'b1000000000110011;
        \commands [403] = 'b1000000010110011;
        \commands [404] = 'b1000000000110011;
        \commands [405] = 'b0001010000000000;
        \commands [406] = 'b1001010000000000;
        \commands [407] = 'b1001010000110100;
        \commands [408] = 'b1001010010110100;
        \commands [409] = 'b1001010000110100;
        \commands [410] = 'b0001010000000000;
        \commands [411] = 'b1001010000000000;
        \commands [412] = 'b1011001000111101;
        \commands [413] = 'b1011001010111101;
        \commands [414] = 'b1011001000111101;
        \commands [415] = 'b0011110100000000;
        \commands [416] = 'b1011110100000000;
        \commands [417] = 'b1011110100111101;
        \commands [418] = 'b1011110110111101;
        \commands [419] = 'b1011110100111101;
        \commands [420] = 'b0011110100000000;
        \commands [421] = 'b1011110100000000;
        \commands [422] = 'b1011001100111101;
        \commands [423] = 'b1011001110111101;
        \commands [424] = 'b1011001100111101;
        \commands [425] = 'b0011010000000000;
        \commands [426] = 'b1011010000000000;
        \commands [427] = 'b1011001000111110;
        \commands [428] = 'b1011001010111110;
        \commands [429] = 'b1011001000111110;
        \commands [430] = 'b0011111000000000;
        \commands [431] = 'b1011111000000000;
        \commands [432] = 'b1011111000111110;
        \commands [433] = 'b1011111010111110;
        \commands [434] = 'b1011111000111110;
        \commands [435] = 'b0011111000000000;
        \commands [436] = 'b1011111000000000;
        \commands [437] = 'b1000000000111110;
        \commands [438] = 'b1000000010111110;
        \commands [439] = 'b1000000000111110;
        \commands [440] = 'b0001010000000000;
        \commands [441] = 'b1001010000000000;
        \commands [442] = 'b1000110100111111;
        \commands [443] = 'b1000110110111111;
        \commands [444] = 'b1000110100111111;
        \commands [445] = 'b0011111100000000;
        \commands [446] = 'b1011111100000000;
        \commands [447] = 'b1011111100111111;
        \commands [448] = 'b1011111110111111;
        \commands [449] = 'b1011111100111111;
        \commands [450] = 'b0011111100000000;
        \commands [451] = 'b1011111100000000;
        \commands [452] = 'b1000000000111111;
        \commands [453] = 'b1000000010111111;
        \commands [454] = 'b1000000000111111;
        \commands [455] = 'b0011010000000000;
        \commands [456] = 'b1011010000000000;
        \commands [457] = 'b1000110101000000;
        \commands [458] = 'b1000110111000000;
        \commands [459] = 'b1000110101000000;
        \commands [460] = 'b0100000000000000;
        \commands [461] = 'b1100000000000000;
        \commands [462] = 'b1100000001000000;
        \commands [463] = 'b1100000011000000;
        \commands [464] = 'b1100000001000000;
        \commands [465] = 'b0100000000000000;
        \commands [466] = 'b1100000000000000;
        \commands [467] = 'b1011001101000000;
        \commands [468] = 'b1011001111000000;
        \commands [469] = 'b1011001101000000;
        \commands [470] = 'b0011110100000000;
        \commands [471] = 'b1011110100000000;
        \commands [472] = 'b1011111001111111;
        \commands [473] = 'b1011111011111111;
        \commands [474] = 'b1011111001111111;
        \commands [475] = 'b0111111100000000;
        \commands [476] = 'b1111111100000000;
        \commands [477] = 'b1111111101111111;
        \commands [478] = 'b1111111111111111;
        \commands [479] = 'b1111111101111111;
        \commands [480] = 'b0011111100000000;
        \commands [481] = 'b1011111100000000;
        \commands [482] = 'b1100000000100001;
        \commands [483] = 'b1100000010100001;
        \commands [484] = 'b1100000000100001;
        \commands [485] = 'b0010000100000000;
        \commands [486] = 'b1010000100000000;
        \commands [487] = 'b1010000100100001;
        \commands [488] = 'b1010000110100001;
        \commands [489] = 'b1010000100100001;
        \commands [490] = 'b0010000100000000;
        \commands [491] = 'b1010000100000000;
        \commands [492] = 'b1111111100100001;
        \commands [493] = 'b1111111110100001;
        \commands [494] = 'b1111111100100001;
        \commands [495] = 'b0000110100000000;
        \commands [496] = 'b1000110100000000;
        \commands [497] = 'b1000000000111101;
        \commands [498] = 'b1000000010111101;
        \commands [499] = 'b1000000000111101;
        \commands [500] = 'b0001010000000000;
        \commands [501] = 'b1001010000000000;
        \commands [502] = 'b1000110100111110;
        \commands [503] = 'b1000110110111110;
        \commands [504] = 'b1000110100111110;
        \commands [505] = 'b0001010000000000;
        \commands [506] = 'b1001010000000000;
        \commands [507] = 'b1000000000111111;
        \commands [508] = 'b1000000010111111;
        \commands [509] = 'b1000000000111111;
        \commands [510] = 'b0011110100000000;
        \commands [511] = 'b1011110100000000;
        \commands [512] = 'b1011111000010100;
        \commands [513] = 'b1011111010010100;
        \commands [514] = 'b1011111000010100;
        \commands [515] = 'b0001010000000000;
        \commands [516] = 'b1001010000000000;
        \commands [517] = 'b1001010000010100;
        \commands [518] = 'b1001010010010100;
        \commands [519] = 'b1001010000010100;
        \commands [520] = 'b0001010000000000;
        \commands [521] = 'b1001010000000000;
        \commands [522] = 'b1011111100010100;
        \commands [523] = 'b1011111110010100;
        \commands [524] = 'b1011111100010100;
        \commands [525] = 'b0000111000000000;
        \commands [526] = 'b1000111000000000;
        \commands [527] = 'b1000111000110010;
        \commands [528] = 'b1000111010110010;
        \commands [529] = 'b1000111000110010;
        \commands [530] = 'b0000000000000000;
        \commands [531] = 'b1000000000000000;
        \commands [532] = 'b1000000000110011;
        \commands [533] = 'b1000000010110011;
        \commands [534] = 'b1000000000110011;
        \commands [535] = 'b0001010000000000;
        \commands [536] = 'b1001010000000000;
        \commands [537] = 'b1001010000110100;
        \commands [538] = 'b1001010010110100;
        \commands [539] = 'b1001010000110100;
        \commands [540] = 'b0001010000000000;
        \commands [541] = 'b1001010000000000;
        \commands [542] = 'b1011001000111101;
        \commands [543] = 'b1011001010111101;
        \commands [544] = 'b1011001000111101;
        \commands [545] = 'b0011110100000000;
        \commands [546] = 'b1011110100000000;
        \commands [547] = 'b1011110100111101;
        \commands [548] = 'b1011110110111101;
        \commands [549] = 'b1011110100111101;
        \commands [550] = 'b0011110100000000;
        \commands [551] = 'b1011110100000000;
        \commands [552] = 'b1011001100111101;
        \commands [553] = 'b1011001110111101;
        \commands [554] = 'b1011001100111101;
        \commands [555] = 'b0011010000000000;
        \commands [556] = 'b1011010000000000;
        \commands [557] = 'b1011001000111110;
        \commands [558] = 'b1011001010111110;
        \commands [559] = 'b1011001000111110;
        \commands [560] = 'b0011111000000000;
        \commands [561] = 'b1011111000000000;
        \commands [562] = 'b1011111000111110;
        \commands [563] = 'b1011111010111110;
        \commands [564] = 'b1011111000111110;
        \commands [565] = 'b0011111000000000;
        \commands [566] = 'b1011111000000000;
        \commands [567] = 'b1000000000111110;
        \commands [568] = 'b1000000010111110;
        \commands [569] = 'b1000000000111110;
        \commands [570] = 'b0001010000000000;
        \commands [571] = 'b1001010000000000;
        \commands [572] = 'b1000111000111111;
        \commands [573] = 'b1000111010111111;
        \commands [574] = 'b1000111000111111;
        \commands [575] = 'b0011111100000000;
        \commands [576] = 'b1011111100000000;
        \commands [577] = 'b1011111100111111;
        \commands [578] = 'b1011111110111111;
        \commands [579] = 'b1011111100111111;
        \commands [580] = 'b0011111100000000;
        \commands [581] = 'b1011111100000000;
        \commands [582] = 'b1000000000111111;
        \commands [583] = 'b1000000010111111;
        \commands [584] = 'b1000000000111111;
        \commands [585] = 'b0011010000000000;
        \commands [586] = 'b1011010000000000;
        \commands [587] = 'b1000111001000000;
        \commands [588] = 'b1000111011000000;
        \commands [589] = 'b1000111001000000;
        \commands [590] = 'b0100000000000000;
        \commands [591] = 'b1100000000000000;
        \commands [592] = 'b1100000001000000;
        \commands [593] = 'b1100000011000000;
        \commands [594] = 'b1100000001000000;
        \commands [595] = 'b0100000000000000;
        \commands [596] = 'b1100000000000000;
        \commands [597] = 'b1011001101000000;
        \commands [598] = 'b1011001111000000;
        \commands [599] = 'b1011001101000000;
        \commands [600] = 'b0011110100000000;
        \commands [601] = 'b1011110100000000;
        \commands [602] = 'b1011111001111111;
        \commands [603] = 'b1011111011111111;
        \commands [604] = 'b1011111001111111;
        \commands [605] = 'b0111111100000000;
        \commands [606] = 'b1111111100000000;
        \commands [607] = 'b1111111101111111;
        \commands [608] = 'b1111111111111111;
        \commands [609] = 'b1111111101111111;
        \commands [610] = 'b0011111100000000;
        \commands [611] = 'b1011111100000000;
        \commands [612] = 'b1100000000100010;
        \commands [613] = 'b1100000010100010;
        \commands [614] = 'b1100000000100010;
        \commands [615] = 'b0010001000000000;
        \commands [616] = 'b1010001000000000;
        \commands [617] = 'b1010001000100010;
        \commands [618] = 'b1010001010100010;
        \commands [619] = 'b1010001000100010;
        \commands [620] = 'b0010001000000000;
        \commands [621] = 'b1010001000000000;
        \commands [622] = 'b1111111100100010;
        \commands [623] = 'b1111111110100010;
        \commands [624] = 'b1111111100100010;
        \commands [625] = 'b0000111000000000;
        \commands [626] = 'b1000111000000000;
        \commands [627] = 'b1000000000111101;
        \commands [628] = 'b1000000010111101;
        \commands [629] = 'b1000000000111101;
        \commands [630] = 'b0001010000000000;
        \commands [631] = 'b1001010000000000;
        \commands [632] = 'b1000111000111110;
        \commands [633] = 'b1000111010111110;
        \commands [634] = 'b1000111000111110;
        \commands [635] = 'b0001010000000000;
        \commands [636] = 'b1001010000000000;
        \commands [637] = 'b1000000000111111;
        \commands [638] = 'b1000000010111111;
        \commands [639] = 'b1000000000111111;
        \commands [640] = 'b0011110100000000;
        \commands [641] = 'b1011110100000000;
        \commands [642] = 'b1011111000010100;
        \commands [643] = 'b1011111010010100;
        \commands [644] = 'b1011111000010100;
        \commands [645] = 'b0001010000000000;
        \commands [646] = 'b1001010000000000;
        \commands [647] = 'b1001010000010100;
        \commands [648] = 'b1001010010010100;
        \commands [649] = 'b1001010000010100;
        \commands [650] = 'b0001010000000000;
        \commands [651] = 'b1001010000000000;
        \commands [652] = 'b1011111100010100;
        \commands [653] = 'b1011111110010100;
        \commands [654] = 'b1011111100010100;
        \commands [655] = 'b0000111100000000;
        \commands [656] = 'b1000111100000000;
        \commands [657] = 'b1000111100110010;
        \commands [658] = 'b1000111110110010;
        \commands [659] = 'b1000111100110010;
        \commands [660] = 'b0000000000000000;
        \commands [661] = 'b1000000000000000;
        \commands [662] = 'b1000000000110011;
        \commands [663] = 'b1000000010110011;
        \commands [664] = 'b1000000000110011;
        \commands [665] = 'b0001010000000000;
        \commands [666] = 'b1001010000000000;
        \commands [667] = 'b1001010000110100;
        \commands [668] = 'b1001010010110100;
        \commands [669] = 'b1001010000110100;
        \commands [670] = 'b0001010000000000;
        \commands [671] = 'b1001010000000000;
        \commands [672] = 'b1011001000111101;
        \commands [673] = 'b1011001010111101;
        \commands [674] = 'b1011001000111101;
        \commands [675] = 'b0011110100000000;
        \commands [676] = 'b1011110100000000;
        \commands [677] = 'b1011110100111101;
        \commands [678] = 'b1011110110111101;
        \commands [679] = 'b1011110100111101;
        \commands [680] = 'b0011110100000000;
        \commands [681] = 'b1011110100000000;
        \commands [682] = 'b1011001100111101;
        \commands [683] = 'b1011001110111101;
        \commands [684] = 'b1011001100111101;
        \commands [685] = 'b0011010000000000;
        \commands [686] = 'b1011010000000000;
        \commands [687] = 'b1011001000111110;
        \commands [688] = 'b1011001010111110;
        \commands [689] = 'b1011001000111110;
        \commands [690] = 'b0011111000000000;
        \commands [691] = 'b1011111000000000;
        \commands [692] = 'b1011111000111110;
        \commands [693] = 'b1011111010111110;
        \commands [694] = 'b1011111000111110;
        \commands [695] = 'b0011111000000000;
        \commands [696] = 'b1011111000000000;
        \commands [697] = 'b1000000000111110;
        \commands [698] = 'b1000000010111110;
        \commands [699] = 'b1000000000111110;
        \commands [700] = 'b0001010000000000;
        \commands [701] = 'b1001010000000000;
        \commands [702] = 'b1000111100111111;
        \commands [703] = 'b1000111110111111;
        \commands [704] = 'b1000111100111111;
        \commands [705] = 'b0011111100000000;
        \commands [706] = 'b1011111100000000;
        \commands [707] = 'b1011111100111111;
        \commands [708] = 'b1011111110111111;
        \commands [709] = 'b1011111100111111;
        \commands [710] = 'b0011111100000000;
        \commands [711] = 'b1011111100000000;
        \commands [712] = 'b1000000000111111;
        \commands [713] = 'b1000000010111111;
        \commands [714] = 'b1000000000111111;
        \commands [715] = 'b0011010000000000;
        \commands [716] = 'b1011010000000000;
        \commands [717] = 'b1000111101000000;
        \commands [718] = 'b1000111111000000;
        \commands [719] = 'b1000111101000000;
        \commands [720] = 'b0100000000000000;
        \commands [721] = 'b1100000000000000;
        \commands [722] = 'b1100000001000000;
        \commands [723] = 'b1100000011000000;
        \commands [724] = 'b1100000001000000;
        \commands [725] = 'b0100000000000000;
        \commands [726] = 'b1100000000000000;
        \commands [727] = 'b1011001101000000;
        \commands [728] = 'b1011001111000000;
        \commands [729] = 'b1011001101000000;
        \commands [730] = 'b0011110100000000;
        \commands [731] = 'b1011110100000000;
        \commands [732] = 'b1011111001111111;
        \commands [733] = 'b1011111011111111;
        \commands [734] = 'b1011111001111111;
        \commands [735] = 'b0111111100000000;
        \commands [736] = 'b1111111100000000;
        \commands [737] = 'b1111111101111111;
        \commands [738] = 'b1111111111111111;
        \commands [739] = 'b1111111101111111;
        \commands [740] = 'b0011111100000000;
        \commands [741] = 'b1011111100000000;
        \commands [742] = 'b1100000000100011;
        \commands [743] = 'b1100000010100011;
        \commands [744] = 'b1100000000100011;
        \commands [745] = 'b0010001100000000;
        \commands [746] = 'b1010001100000000;
        \commands [747] = 'b1010001100100011;
        \commands [748] = 'b1010001110100011;
        \commands [749] = 'b1010001100100011;
        \commands [750] = 'b0010001100000000;
        \commands [751] = 'b1010001100000000;
        \commands [752] = 'b1111111100100011;
        \commands [753] = 'b1111111110100011;
        \commands [754] = 'b1111111100100011;
        \commands [755] = 'b0000111100000000;
        \commands [756] = 'b1000111100000000;
        \commands [757] = 'b1000000000111101;
        \commands [758] = 'b1000000010111101;
        \commands [759] = 'b1000000000111101;
        \commands [760] = 'b0001010000000000;
        \commands [761] = 'b1001010000000000;
        \commands [762] = 'b1000111100111110;
        \commands [763] = 'b1000111110111110;
        \commands [764] = 'b1000111100111110;
        \commands [765] = 'b0001010000000000;
        \commands [766] = 'b1001010000000000;
        \commands [767] = 'b1000000000111111;
        \commands [768] = 'b1000000010111111;
        \commands [769] = 'b1000000000111111;
        \commands [770] = 'b0011110100000000;
        \commands [771] = 'b1011110100000000;
        \commands [772] = 'b1011111000010100;
        \commands [773] = 'b1011111010010100;
        \commands [774] = 'b1011111000010100;
        \commands [775] = 'b0001010000000000;
        \commands [776] = 'b1001010000000000;
        \commands [777] = 'b1001010000010100;
        \commands [778] = 'b1001010010010100;
        \commands [779] = 'b1001010000010100;
        \commands [780] = 'b0001010000000000;
        \commands [781] = 'b1001010000000000;
        \commands [782] = 'b1011111100010100;
        \commands [783] = 'b1011111110010100;
        \commands [784] = 'b1011111100010100;
        \commands [785] = 'b0001000000000000;
        \commands [786] = 'b1001000000000000;
        \commands [787] = 'b1001000000110010;
        \commands [788] = 'b1001000010110010;
        \commands [789] = 'b1001000000110010;
        \commands [790] = 'b0000000000000000;
        \commands [791] = 'b1000000000000000;
        \commands [792] = 'b1000000000110011;
        \commands [793] = 'b1000000010110011;
        \commands [794] = 'b1000000000110011;
        \commands [795] = 'b0001010000000000;
        \commands [796] = 'b1001010000000000;
        \commands [797] = 'b1001010000110100;
        \commands [798] = 'b1001010010110100;
        \commands [799] = 'b1001010000110100;
        \commands [800] = 'b0001010000000000;
        \commands [801] = 'b1001010000000000;
        \commands [802] = 'b1011001000111101;
        \commands [803] = 'b1011001010111101;
        \commands [804] = 'b1011001000111101;
        \commands [805] = 'b0011110100000000;
        \commands [806] = 'b1011110100000000;
        \commands [807] = 'b1011110100111101;
        \commands [808] = 'b1011110110111101;
        \commands [809] = 'b1011110100111101;
        \commands [810] = 'b0011110100000000;
        \commands [811] = 'b1011110100000000;
        \commands [812] = 'b1011001100111101;
        \commands [813] = 'b1011001110111101;
        \commands [814] = 'b1011001100111101;
        \commands [815] = 'b0011010000000000;
        \commands [816] = 'b1011010000000000;
        \commands [817] = 'b1011001000111110;
        \commands [818] = 'b1011001010111110;
        \commands [819] = 'b1011001000111110;
        \commands [820] = 'b0011111000000000;
        \commands [821] = 'b1011111000000000;
        \commands [822] = 'b1011111000111110;
        \commands [823] = 'b1011111010111110;
        \commands [824] = 'b1011111000111110;
        \commands [825] = 'b0011111000000000;
        \commands [826] = 'b1011111000000000;
        \commands [827] = 'b1000000000111110;
        \commands [828] = 'b1000000010111110;
        \commands [829] = 'b1000000000111110;
        \commands [830] = 'b0001010000000000;
        \commands [831] = 'b1001010000000000;
        \commands [832] = 'b1001000000111111;
        \commands [833] = 'b1001000010111111;
        \commands [834] = 'b1001000000111111;
        \commands [835] = 'b0011111100000000;
        \commands [836] = 'b1011111100000000;
        \commands [837] = 'b1011111100111111;
        \commands [838] = 'b1011111110111111;
        \commands [839] = 'b1011111100111111;
        \commands [840] = 'b0011111100000000;
        \commands [841] = 'b1011111100000000;
        \commands [842] = 'b1000000000111111;
        \commands [843] = 'b1000000010111111;
        \commands [844] = 'b1000000000111111;
        \commands [845] = 'b0011010000000000;
        \commands [846] = 'b1011010000000000;
        \commands [847] = 'b1001000001000000;
        \commands [848] = 'b1001000011000000;
        \commands [849] = 'b1001000001000000;
        \commands [850] = 'b0100000000000000;
        \commands [851] = 'b1100000000000000;
        \commands [852] = 'b1100000001000000;
        \commands [853] = 'b1100000011000000;
        \commands [854] = 'b1100000001000000;
        \commands [855] = 'b0100000000000000;
        \commands [856] = 'b1100000000000000;
        \commands [857] = 'b1011001101000000;
        \commands [858] = 'b1011001111000000;
        \commands [859] = 'b1011001101000000;
        \commands [860] = 'b0011110100000000;
        \commands [861] = 'b1011110100000000;
        \commands [862] = 'b1011111001111111;
        \commands [863] = 'b1011111011111111;
        \commands [864] = 'b1011111001111111;
        \commands [865] = 'b0111111100000000;
        \commands [866] = 'b1111111100000000;
        \commands [867] = 'b1111111101111111;
        \commands [868] = 'b1111111111111111;
        \commands [869] = 'b1111111101111111;
        \commands [870] = 'b0011111100000000;
        \commands [871] = 'b1011111100000000;
        \commands [872] = 'b1100000000100100;
        \commands [873] = 'b1100000010100100;
        \commands [874] = 'b1100000000100100;
        \commands [875] = 'b0010010000000000;
        \commands [876] = 'b1010010000000000;
        \commands [877] = 'b1010010000100100;
        \commands [878] = 'b1010010010100100;
        \commands [879] = 'b1010010000100100;
        \commands [880] = 'b0010010000000000;
        \commands [881] = 'b1010010000000000;
        \commands [882] = 'b1111111100100100;
        \commands [883] = 'b1111111110100100;
        \commands [884] = 'b1111111100100100;
        \commands [885] = 'b0001000000000000;
        \commands [886] = 'b1001000000000000;
        \commands [887] = 'b1000000000111101;
        \commands [888] = 'b1000000010111101;
        \commands [889] = 'b1000000000111101;
        \commands [890] = 'b0001010000000000;
        \commands [891] = 'b1001010000000000;
        \commands [892] = 'b1001000000111110;
        \commands [893] = 'b1001000010111110;
        \commands [894] = 'b1001000000111110;
        \commands [895] = 'b0001010000000000;
        \commands [896] = 'b1001010000000000;
        \commands [897] = 'b1000000000111111;
        \commands [898] = 'b1000000010111111;
        \commands [899] = 'b1000000000111111;
        \commands [900] = 'b0011110100000000;
        \commands [901] = 'b1011110100000000;
        \commands [902] = 'b1011111000010100;
        \commands [903] = 'b1011111010010100;
        \commands [904] = 'b1011111000010100;
        \commands [905] = 'b0001010000000000;
        \commands [906] = 'b1001010000000000;
        \commands [907] = 'b1001010000010100;
        \commands [908] = 'b1001010010010100;
        \commands [909] = 'b1001010000010100;
        \commands [910] = 'b0001010000000000;
        \commands [911] = 'b1001010000000000;
        \commands [912] = 'b1011111100010100;
        \commands [913] = 'b1011111110010100;
        \commands [914] = 'b1011111100010100;
        \commands [915] = 'b0001000100000000;
        \commands [916] = 'b1001000100000000;
        \commands [917] = 'b1001000100110010;
        \commands [918] = 'b1001000110110010;
        \commands [919] = 'b1001000100110010;
        \commands [920] = 'b0000000000000000;
        \commands [921] = 'b1000000000000000;
        \commands [922] = 'b1000000000110011;
        \commands [923] = 'b1000000010110011;
        \commands [924] = 'b1000000000110011;
        \commands [925] = 'b0001010000000000;
        \commands [926] = 'b1001010000000000;
        \commands [927] = 'b1001010000110100;
        \commands [928] = 'b1001010010110100;
        \commands [929] = 'b1001010000110100;
        \commands [930] = 'b0001010000000000;
        \commands [931] = 'b1001010000000000;
        \commands [932] = 'b1011001000111101;
        \commands [933] = 'b1011001010111101;
        \commands [934] = 'b1011001000111101;
        \commands [935] = 'b0011110100000000;
        \commands [936] = 'b1011110100000000;
        \commands [937] = 'b1011110100111101;
        \commands [938] = 'b1011110110111101;
        \commands [939] = 'b1011110100111101;
        \commands [940] = 'b0011110100000000;
        \commands [941] = 'b1011110100000000;
        \commands [942] = 'b1011001100111101;
        \commands [943] = 'b1011001110111101;
        \commands [944] = 'b1011001100111101;
        \commands [945] = 'b0011010000000000;
        \commands [946] = 'b1011010000000000;
        \commands [947] = 'b1011001000111110;
        \commands [948] = 'b1011001010111110;
        \commands [949] = 'b1011001000111110;
        \commands [950] = 'b0011111000000000;
        \commands [951] = 'b1011111000000000;
        \commands [952] = 'b1011111000111110;
        \commands [953] = 'b1011111010111110;
        \commands [954] = 'b1011111000111110;
        \commands [955] = 'b0011111000000000;
        \commands [956] = 'b1011111000000000;
        \commands [957] = 'b1000000000111110;
        \commands [958] = 'b1000000010111110;
        \commands [959] = 'b1000000000111110;
        \commands [960] = 'b0001010000000000;
        \commands [961] = 'b1001010000000000;
        \commands [962] = 'b1001000100111111;
        \commands [963] = 'b1001000110111111;
        \commands [964] = 'b1001000100111111;
        \commands [965] = 'b0011111100000000;
        \commands [966] = 'b1011111100000000;
        \commands [967] = 'b1011111100111111;
        \commands [968] = 'b1011111110111111;
        \commands [969] = 'b1011111100111111;
        \commands [970] = 'b0011111100000000;
        \commands [971] = 'b1011111100000000;
        \commands [972] = 'b1000000000111111;
        \commands [973] = 'b1000000010111111;
        \commands [974] = 'b1000000000111111;
        \commands [975] = 'b0011010000000000;
        \commands [976] = 'b1011010000000000;
        \commands [977] = 'b1001000101000000;
        \commands [978] = 'b1001000111000000;
        \commands [979] = 'b1001000101000000;
        \commands [980] = 'b0100000000000000;
        \commands [981] = 'b1100000000000000;
        \commands [982] = 'b1100000001000000;
        \commands [983] = 'b1100000011000000;
        \commands [984] = 'b1100000001000000;
        \commands [985] = 'b0100000000000000;
        \commands [986] = 'b1100000000000000;
        \commands [987] = 'b1011001101000000;
        \commands [988] = 'b1011001111000000;
        \commands [989] = 'b1011001101000000;
        \commands [990] = 'b0011110100000000;
        \commands [991] = 'b1011110100000000;
        \commands [992] = 'b1011111001111111;
        \commands [993] = 'b1011111011111111;
        \commands [994] = 'b1011111001111111;
        \commands [995] = 'b0111111100000000;
        \commands [996] = 'b1111111100000000;
        \commands [997] = 'b1111111101111111;
        \commands [998] = 'b1111111111111111;
        \commands [999] = 'b1111111101111111;
        \commands [1000] = 'b0011111100000000;
        \commands [1001] = 'b1011111100000000;
        \commands [1002] = 'b1100000000100101;
        \commands [1003] = 'b1100000010100101;
        \commands [1004] = 'b1100000000100101;
        \commands [1005] = 'b0010010100000000;
        \commands [1006] = 'b1010010100000000;
        \commands [1007] = 'b1010010100100101;
        \commands [1008] = 'b1010010110100101;
        \commands [1009] = 'b1010010100100101;
        \commands [1010] = 'b0010010100000000;
        \commands [1011] = 'b1010010100000000;
        \commands [1012] = 'b1111111100100101;
        \commands [1013] = 'b1111111110100101;
        \commands [1014] = 'b1111111100100101;
        \commands [1015] = 'b0001000100000000;
        \commands [1016] = 'b1001000100000000;
        \commands [1017] = 'b1000000000111101;
        \commands [1018] = 'b1000000010111101;
        \commands [1019] = 'b1000000000111101;
        \commands [1020] = 'b0001010000000000;
        \commands [1021] = 'b1001010000000000;
        \commands [1022] = 'b1001000100111110;
        \commands [1023] = 'b1001000110111110;
        \commands [1024] = 'b1001000100111110;
        \commands [1025] = 'b0001010000000000;
        \commands [1026] = 'b1001010000000000;
        \commands [1027] = 'b1000000000111111;
        \commands [1028] = 'b1000000010111111;
        \commands [1029] = 'b1000000000111111;
        \commands [1030] = 'b0011110100000000;
        \commands [1031] = 'b1011110100000000;
        \commands [1032] = 'b1011111000010100;
        \commands [1033] = 'b1011111010010100;
        \commands [1034] = 'b1011111000010100;
        \commands [1035] = 'b0001010000000000;
        \commands [1036] = 'b1001010000000000;
        \commands [1037] = 'b1001010000010100;
        \commands [1038] = 'b1001010010010100;
        \commands [1039] = 'b1001010000010100;
        \commands [1040] = 'b0001010000000000;
        \commands [1041] = 'b1001010000000000;
        \commands [1042] = 'b1011111100010100;
        \commands [1043] = 'b1011111110010100;
        \commands [1044] = 'b1011111100010100;
        \commands [1045] = 'b0001111000000000;
        \commands [1046] = 'b1001111000000000;
        \commands [1047] = 'b1001111000001010;
        \commands [1048] = 'b1001111010001010;
        \commands [1049] = 'b1001111000001010;
        \commands [1050] = 'b0000101000000001;
        \commands [1051] = 'b1000101000000001;
        \commands [1052] = 'b1000101000001010;
        \commands [1053] = 'b1000101010001010;
        \commands [1054] = 'b1000101000001010;
        \commands [1055] = 'b0001111100000000;
        \commands [1056] = 'b1001111100000000;
        \commands [1057] = 'b1001111100001011;
        \commands [1058] = 'b1001111110001011;
        \commands [1059] = 'b1001111100001011;
        \commands [1060] = 'b0000101100000001;
        \commands [1061] = 'b1000101100000001;
        \commands [1062] = 'b1000101100001011;
        \commands [1063] = 'b1000101110001011;
        \commands [1064] = 'b1000101100001011;
        \commands [1065] = 'b0010000000000000;
        \commands [1066] = 'b1010000000000000;
        \commands [1067] = 'b1010000000001100;
        \commands [1068] = 'b1010000010001100;
        \commands [1069] = 'b1010000000001100;
        \commands [1070] = 'b0000110000000001;
        \commands [1071] = 'b1000110000000001;
        \commands [1072] = 'b1000110000001100;
        \commands [1073] = 'b1000110010001100;
        \commands [1074] = 'b1000110000001100;
        \commands [1075] = 'b0010000100000000;
        \commands [1076] = 'b1010000100000000;
        \commands [1077] = 'b1010000100001101;
        \commands [1078] = 'b1010000110001101;
        \commands [1079] = 'b1010000100001101;
        \commands [1080] = 'b0000110100000001;
        \commands [1081] = 'b1000110100000001;
        \commands [1082] = 'b1000110100001101;
        \commands [1083] = 'b1000110110001101;
        \commands [1084] = 'b1000110100001101;
        \commands [1085] = 'b0010001000000000;
        \commands [1086] = 'b1010001000000000;
        \commands [1087] = 'b1010001000001110;
        \commands [1088] = 'b1010001010001110;
        \commands [1089] = 'b1010001000001110;
        \commands [1090] = 'b0000111000000001;
        \commands [1091] = 'b1000111000000001;
        \commands [1092] = 'b1000111000001110;
        \commands [1093] = 'b1000111010001110;
        \commands [1094] = 'b1000111000001110;
        \commands [1095] = 'b0010001100000000;
        \commands [1096] = 'b1010001100000000;
        \commands [1097] = 'b1010001100001111;
        \commands [1098] = 'b1010001110001111;
        \commands [1099] = 'b1010001100001111;
        \commands [1100] = 'b0000111100000001;
        \commands [1101] = 'b1000111100000001;
        \commands [1102] = 'b1000111100001111;
        \commands [1103] = 'b1000111110001111;
        \commands [1104] = 'b1000111100001111;
        \commands [1105] = 'b0010010000000000;
        \commands [1106] = 'b1010010000000000;
        \commands [1107] = 'b1010010000010000;
        \commands [1108] = 'b1010010010010000;
        \commands [1109] = 'b1010010000010000;
        \commands [1110] = 'b0001000000000001;
        \commands [1111] = 'b1001000000000001;
        \commands [1112] = 'b1001000000010000;
        \commands [1113] = 'b1001000010010000;
        \commands [1114] = 'b1001000000010000;
        \commands [1115] = 'b0010010100000000;
        \commands [1116] = 'b1010010100000000;
        \commands [1117] = 'b1010010100010001;
        \commands [1118] = 'b1010010110010001;
        \commands [1119] = 'b1010010100010001;
        \commands [1120] = 'b0001000100000001;
        \commands [1121] = 'b1001000100000001;
        \commands [1122] = 'b1001000100010001;
        \commands [1123] = 'b1001000110010001;
        \commands [1124] = 'b1001000100010001;
    end
    always @(posedge \clk ) begin
        
    end
    assign _e_3741 = \read_idx [10:0];
    assign \mem_out  = \commands [_e_3741];
    assign \a  = \s1_mem_out [15:8];
    assign \b  = \s1_mem_out [7:0];
    assign _e_3748 = {\a , \b };
    assign output__ = _e_3748;
endmodule